`include "data/modules/LSmitll_XORT_v2p1_selfcontained.v"
`include "data/modules/LSmitll_AND2T_v2p1_selfcontained.v"
`include "data/modules/LSmitll_SPLITT_v2p1_selfcontained.v"
`include "data/modules/LSmitll_OR2T_v2p1_selfcontained.v"
`include "data/modules/LSmitll_DFFT_v2p1_selfcontained.v"
`timescale 1ps/100fs
module KSA8 (
	a0,
	b0,
	sum0,
	sum1,
	sum2,
	sum3,
	sum4,
	sum5,
	sum6,
	sum7,
	cout,
	a1,
	a2,
	a3,
	a4,
	a5,
	a6,
	a7,
	b1,
	b2,
	b3,
	b4,
	b5,
	b6,
	b7,
	cin,
	clk
);
input
	a0,b0,a1,a2,a3,a4,a5,a6,a7,b1,b2,b3,b4,b5,b6,b7,cin,clk;

output
	sum0,sum1,sum2,sum3,sum4,sum5,sum6,sum7,cout;

reg  [827:0] net_r = 0;
wire [827:0] net_w;
assign net_w[1] = a0;
assign net_w[9] = b0;
assign net_w[64] = a1;
assign net_w[68] = a2;
assign net_w[74] = a3;
assign net_w[82] = a4;
assign net_w[92] = a5;
assign net_w[104] = a6;
assign net_w[118] = a7;
assign net_w[120] = b1;
assign net_w[124] = b2;
assign net_w[130] = b3;
assign net_w[138] = b4;
assign net_w[148] = b5;
assign net_w[160] = b6;
assign net_w[174] = b7;
assign net_w[175] = cin;
assign net_w[332] = clk;
assign sum0 = net_r[54];
assign sum1 = net_r[55];
assign sum2 = net_r[56];
assign sum3 = net_r[57];
assign sum4 = net_r[58];
assign sum5 = net_r[59];
assign sum6 = net_r[60];
assign sum7 = net_r[61];
assign cout = net_r[62];
always @(posedge net_w[1] or negedge net_w[1]) begin
	#1.47213 net_r[1] <= net_w[1];
end
always @(posedge net_w[2] or negedge net_w[2]) begin
	#0.84122 net_r[2] <= net_w[2];
end
always @(posedge net_w[3] or negedge net_w[3]) begin
	#1.78759 net_r[3] <= net_w[3];
end
always @(posedge net_w[4] or negedge net_w[4]) begin
	#0.42061 net_r[4] <= net_w[4];
end
always @(posedge net_w[5] or negedge net_w[5]) begin
	#1.9979 net_r[5] <= net_w[5];
end
always @(posedge net_w[6] or negedge net_w[6]) begin
	#1.68244 net_r[6] <= net_w[6];
end
always @(posedge net_w[7] or negedge net_w[7]) begin
	#3.04942 net_r[7] <= net_w[7];
end
always @(posedge net_w[8] or negedge net_w[8]) begin
	#2.52366 net_r[8] <= net_w[8];
end
always @(posedge net_w[9] or negedge net_w[9]) begin
	#1.26183 net_r[9] <= net_w[9];
end
always @(posedge net_w[10] or negedge net_w[10]) begin
	#0.630915 net_r[10] <= net_w[10];
end
always @(posedge net_w[11] or negedge net_w[11]) begin
	#1.36698 net_r[11] <= net_w[11];
end
always @(posedge net_w[12] or negedge net_w[12]) begin
	#0.736067 net_r[12] <= net_w[12];
end
always @(posedge net_w[13] or negedge net_w[13]) begin
	#0.736067 net_r[13] <= net_w[13];
end
always @(posedge net_w[14] or negedge net_w[14]) begin
	#0.84122 net_r[14] <= net_w[14];
end
always @(posedge net_w[15] or negedge net_w[15]) begin
	#0.42061 net_r[15] <= net_w[15];
end
always @(posedge net_w[16] or negedge net_w[16]) begin
	#0.736067 net_r[16] <= net_w[16];
end
always @(posedge net_w[17] or negedge net_w[17]) begin
	#1.36698 net_r[17] <= net_w[17];
end
always @(posedge net_w[18] or negedge net_w[18]) begin
	#0.42061 net_r[18] <= net_w[18];
end
always @(posedge net_w[19] or negedge net_w[19]) begin
	#3.57518 net_r[19] <= net_w[19];
end
always @(posedge net_w[20] or negedge net_w[20]) begin
	#1.68244 net_r[20] <= net_w[20];
end
always @(posedge net_w[21] or negedge net_w[21]) begin
	#1.47213 net_r[21] <= net_w[21];
end
always @(posedge net_w[22] or negedge net_w[22]) begin
	#1.57729 net_r[22] <= net_w[22];
end
always @(posedge net_w[23] or negedge net_w[23]) begin
	#0.84122 net_r[23] <= net_w[23];
end
always @(posedge net_w[24] or negedge net_w[24]) begin
	#5.67823 net_r[24] <= net_w[24];
end
always @(posedge net_w[25] or negedge net_w[25]) begin
	#2.10305 net_r[25] <= net_w[25];
end
always @(posedge net_w[26] or negedge net_w[26]) begin
	#1.05152 net_r[26] <= net_w[26];
end
always @(posedge net_w[27] or negedge net_w[27]) begin
	#6.51945 net_r[27] <= net_w[27];
end
always @(posedge net_w[28] or negedge net_w[28]) begin
	#0.946372 net_r[28] <= net_w[28];
end
always @(posedge net_w[29] or negedge net_w[29]) begin
	#1.57729 net_r[29] <= net_w[29];
end
always @(posedge net_w[30] or negedge net_w[30]) begin
	#5.25762 net_r[30] <= net_w[30];
end
always @(posedge net_w[31] or negedge net_w[31]) begin
	#7.67613 net_r[31] <= net_w[31];
end
always @(posedge net_w[32] or negedge net_w[32]) begin
	#5.46793 net_r[32] <= net_w[32];
end
always @(posedge net_w[33] or negedge net_w[33]) begin
	#5.78339 net_r[33] <= net_w[33];
end
always @(posedge net_w[34] or negedge net_w[34]) begin
	#2.2082 net_r[34] <= net_w[34];
end
always @(posedge net_w[35] or negedge net_w[35]) begin
	#1.26183 net_r[35] <= net_w[35];
end
always @(posedge net_w[36] or negedge net_w[36]) begin
	#10.4101 net_r[36] <= net_w[36];
end
always @(posedge net_w[37] or negedge net_w[37]) begin
	#9.04311 net_r[37] <= net_w[37];
end
always @(posedge net_w[38] or negedge net_w[38]) begin
	#7.99159 net_r[38] <= net_w[38];
end
always @(posedge net_w[39] or negedge net_w[39]) begin
	#1.05152 net_r[39] <= net_w[39];
end
always @(posedge net_w[40] or negedge net_w[40]) begin
	#4.2061 net_r[40] <= net_w[40];
end
always @(posedge net_w[41] or negedge net_w[41]) begin
	#9.98948 net_r[41] <= net_w[41];
end
always @(posedge net_w[42] or negedge net_w[42]) begin
	#13.2492 net_r[42] <= net_w[42];
end
always @(posedge net_w[43] or negedge net_w[43]) begin
	#11.8822 net_r[43] <= net_w[43];
end
always @(posedge net_w[44] or negedge net_w[44]) begin
	#2.10305 net_r[44] <= net_w[44];
end
always @(posedge net_w[45] or negedge net_w[45]) begin
	#1.36698 net_r[45] <= net_w[45];
end
always @(posedge net_w[46] or negedge net_w[46]) begin
	#12.3028 net_r[46] <= net_w[46];
end
always @(posedge net_w[47] or negedge net_w[47]) begin
	#9.98948 net_r[47] <= net_w[47];
end
always @(posedge net_w[48] or negedge net_w[48]) begin
	#11.2513 net_r[48] <= net_w[48];
end
always @(posedge net_w[49] or negedge net_w[49]) begin
	#1.78759 net_r[49] <= net_w[49];
end
always @(posedge net_w[50] or negedge net_w[50]) begin
	#2.41851 net_r[50] <= net_w[50];
end
always @(posedge net_w[51] or negedge net_w[51]) begin
	#14.511 net_r[51] <= net_w[51];
end
always @(posedge net_w[52] or negedge net_w[52]) begin
	#11.041 net_r[52] <= net_w[52];
end
always @(posedge net_w[53] or negedge net_w[53]) begin
	#4.2061 net_r[53] <= net_w[53];
end
always @(posedge net_w[54] or negedge net_w[54]) begin
	#10.5152 net_r[54] <= net_w[54];
end
always @(posedge net_w[55] or negedge net_w[55]) begin
	#8.93796 net_r[55] <= net_w[55];
end
always @(posedge net_w[56] or negedge net_w[56]) begin
	#9.88433 net_r[56] <= net_w[56];
end
always @(posedge net_w[57] or negedge net_w[57]) begin
	#9.98948 net_r[57] <= net_w[57];
end
always @(posedge net_w[58] or negedge net_w[58]) begin
	#9.98948 net_r[58] <= net_w[58];
end
always @(posedge net_w[59] or negedge net_w[59]) begin
	#8.72766 net_r[59] <= net_w[59];
end
always @(posedge net_w[60] or negedge net_w[60]) begin
	#7.46583 net_r[60] <= net_w[60];
end
always @(posedge net_w[61] or negedge net_w[61]) begin
	#8.30705 net_r[61] <= net_w[61];
end
always @(posedge net_w[62] or negedge net_w[62]) begin
	#4.10095 net_r[62] <= net_w[62];
end
always @(posedge net_w[63] or negedge net_w[63]) begin
	#2.2082 net_r[63] <= net_w[63];
end
always @(posedge net_w[64] or negedge net_w[64]) begin
	#2.10305 net_r[64] <= net_w[64];
end
always @(posedge net_w[65] or negedge net_w[65]) begin
	#3.04942 net_r[65] <= net_w[65];
end
always @(posedge net_w[66] or negedge net_w[66]) begin
	#1.47213 net_r[66] <= net_w[66];
end
always @(posedge net_w[67] or negedge net_w[67]) begin
	#2.2082 net_r[67] <= net_w[67];
end
always @(posedge net_w[68] or negedge net_w[68]) begin
	#2.10305 net_r[68] <= net_w[68];
end
always @(posedge net_w[69] or negedge net_w[69]) begin
	#1.89274 net_r[69] <= net_w[69];
end
always @(posedge net_w[70] or negedge net_w[70]) begin
	#2.41851 net_r[70] <= net_w[70];
end
always @(posedge net_w[71] or negedge net_w[71]) begin
	#2.94427 net_r[71] <= net_w[71];
end
always @(posedge net_w[72] or negedge net_w[72]) begin
	#1.36698 net_r[72] <= net_w[72];
end
always @(posedge net_w[73] or negedge net_w[73]) begin
	#2.2082 net_r[73] <= net_w[73];
end
always @(posedge net_w[74] or negedge net_w[74]) begin
	#1.9979 net_r[74] <= net_w[74];
end
always @(posedge net_w[75] or negedge net_w[75]) begin
	#3.36488 net_r[75] <= net_w[75];
end
always @(posedge net_w[76] or negedge net_w[76]) begin
	#1.26183 net_r[76] <= net_w[76];
end
always @(posedge net_w[77] or negedge net_w[77]) begin
	#1.9979 net_r[77] <= net_w[77];
end
always @(posedge net_w[78] or negedge net_w[78]) begin
	#2.31335 net_r[78] <= net_w[78];
end
always @(posedge net_w[79] or negedge net_w[79]) begin
	#2.83912 net_r[79] <= net_w[79];
end
always @(posedge net_w[80] or negedge net_w[80]) begin
	#1.26183 net_r[80] <= net_w[80];
end
always @(posedge net_w[81] or negedge net_w[81]) begin
	#2.2082 net_r[81] <= net_w[81];
end
always @(posedge net_w[82] or negedge net_w[82]) begin
	#1.89274 net_r[82] <= net_w[82];
end
always @(posedge net_w[83] or negedge net_w[83]) begin
	#2.73396 net_r[83] <= net_w[83];
end
always @(posedge net_w[84] or negedge net_w[84]) begin
	#2.10305 net_r[84] <= net_w[84];
end
always @(posedge net_w[85] or negedge net_w[85]) begin
	#3.36488 net_r[85] <= net_w[85];
end
always @(posedge net_w[86] or negedge net_w[86]) begin
	#1.15668 net_r[86] <= net_w[86];
end
always @(posedge net_w[87] or negedge net_w[87]) begin
	#1.78759 net_r[87] <= net_w[87];
end
always @(posedge net_w[88] or negedge net_w[88]) begin
	#2.10305 net_r[88] <= net_w[88];
end
always @(posedge net_w[89] or negedge net_w[89]) begin
	#2.73396 net_r[89] <= net_w[89];
end
always @(posedge net_w[90] or negedge net_w[90]) begin
	#1.26183 net_r[90] <= net_w[90];
end
always @(posedge net_w[91] or negedge net_w[91]) begin
	#2.2082 net_r[91] <= net_w[91];
end
always @(posedge net_w[92] or negedge net_w[92]) begin
	#1.89274 net_r[92] <= net_w[92];
end
always @(posedge net_w[93] or negedge net_w[93]) begin
	#4.10095 net_r[93] <= net_w[93];
end
always @(posedge net_w[94] or negedge net_w[94]) begin
	#1.78759 net_r[94] <= net_w[94];
end
always @(posedge net_w[95] or negedge net_w[95]) begin
	#2.73396 net_r[95] <= net_w[95];
end
always @(posedge net_w[96] or negedge net_w[96]) begin
	#2.10305 net_r[96] <= net_w[96];
end
always @(posedge net_w[97] or negedge net_w[97]) begin
	#3.25973 net_r[97] <= net_w[97];
end
always @(posedge net_w[98] or negedge net_w[98]) begin
	#1.15668 net_r[98] <= net_w[98];
end
always @(posedge net_w[99] or negedge net_w[99]) begin
	#1.78759 net_r[99] <= net_w[99];
end
always @(posedge net_w[100] or negedge net_w[100]) begin
	#1.9979 net_r[100] <= net_w[100];
end
always @(posedge net_w[101] or negedge net_w[101]) begin
	#2.62881 net_r[101] <= net_w[101];
end
always @(posedge net_w[102] or negedge net_w[102]) begin
	#1.15668 net_r[102] <= net_w[102];
end
always @(posedge net_w[103] or negedge net_w[103]) begin
	#2.2082 net_r[103] <= net_w[103];
end
always @(posedge net_w[104] or negedge net_w[104]) begin
	#1.78759 net_r[104] <= net_w[104];
end
always @(posedge net_w[105] or negedge net_w[105]) begin
	#3.89064 net_r[105] <= net_w[105];
end
always @(posedge net_w[106] or negedge net_w[106]) begin
	#3.04942 net_r[106] <= net_w[106];
end
always @(posedge net_w[107] or negedge net_w[107]) begin
	#3.78549 net_r[107] <= net_w[107];
end
always @(posedge net_w[108] or negedge net_w[108]) begin
	#1.9979 net_r[108] <= net_w[108];
end
always @(posedge net_w[109] or negedge net_w[109]) begin
	#3.04942 net_r[109] <= net_w[109];
end
always @(posedge net_w[110] or negedge net_w[110]) begin
	#2.10305 net_r[110] <= net_w[110];
end
always @(posedge net_w[111] or negedge net_w[111]) begin
	#3.25973 net_r[111] <= net_w[111];
end
always @(posedge net_w[112] or negedge net_w[112]) begin
	#1.15668 net_r[112] <= net_w[112];
end
always @(posedge net_w[113] or negedge net_w[113]) begin
	#1.89274 net_r[113] <= net_w[113];
end
always @(posedge net_w[114] or negedge net_w[114]) begin
	#1.89274 net_r[114] <= net_w[114];
end
always @(posedge net_w[115] or negedge net_w[115]) begin
	#2.52366 net_r[115] <= net_w[115];
end
always @(posedge net_w[116] or negedge net_w[116]) begin
	#1.05152 net_r[116] <= net_w[116];
end
always @(posedge net_w[117] or negedge net_w[117]) begin
	#2.2082 net_r[117] <= net_w[117];
end
always @(posedge net_w[118] or negedge net_w[118]) begin
	#1.68244 net_r[118] <= net_w[118];
end
always @(posedge net_w[119] or negedge net_w[119]) begin
	#1.9979 net_r[119] <= net_w[119];
end
always @(posedge net_w[120] or negedge net_w[120]) begin
	#1.89274 net_r[120] <= net_w[120];
end
always @(posedge net_w[121] or negedge net_w[121]) begin
	#1.78759 net_r[121] <= net_w[121];
end
always @(posedge net_w[122] or negedge net_w[122]) begin
	#1.26183 net_r[122] <= net_w[122];
end
always @(posedge net_w[123] or negedge net_w[123]) begin
	#1.78759 net_r[123] <= net_w[123];
end
always @(posedge net_w[124] or negedge net_w[124]) begin
	#1.78759 net_r[124] <= net_w[124];
end
always @(posedge net_w[125] or negedge net_w[125]) begin
	#2.41851 net_r[125] <= net_w[125];
end
always @(posedge net_w[126] or negedge net_w[126]) begin
	#1.9979 net_r[126] <= net_w[126];
end
always @(posedge net_w[127] or negedge net_w[127]) begin
	#1.89274 net_r[127] <= net_w[127];
end
always @(posedge net_w[128] or negedge net_w[128]) begin
	#1.15668 net_r[128] <= net_w[128];
end
always @(posedge net_w[129] or negedge net_w[129]) begin
	#1.9979 net_r[129] <= net_w[129];
end
always @(posedge net_w[130] or negedge net_w[130]) begin
	#1.78759 net_r[130] <= net_w[130];
end
always @(posedge net_w[131] or negedge net_w[131]) begin
	#2.41851 net_r[131] <= net_w[131];
end
always @(posedge net_w[132] or negedge net_w[132]) begin
	#1.36698 net_r[132] <= net_w[132];
end
always @(posedge net_w[133] or negedge net_w[133]) begin
	#2.41851 net_r[133] <= net_w[133];
end
always @(posedge net_w[134] or negedge net_w[134]) begin
	#1.78759 net_r[134] <= net_w[134];
end
always @(posedge net_w[135] or negedge net_w[135]) begin
	#1.89274 net_r[135] <= net_w[135];
end
always @(posedge net_w[136] or negedge net_w[136]) begin
	#1.05152 net_r[136] <= net_w[136];
end
always @(posedge net_w[137] or negedge net_w[137]) begin
	#1.78759 net_r[137] <= net_w[137];
end
always @(posedge net_w[138] or negedge net_w[138]) begin
	#1.68244 net_r[138] <= net_w[138];
end
always @(posedge net_w[139] or negedge net_w[139]) begin
	#2.10305 net_r[139] <= net_w[139];
end
always @(posedge net_w[140] or negedge net_w[140]) begin
	#1.47213 net_r[140] <= net_w[140];
end
always @(posedge net_w[141] or negedge net_w[141]) begin
	#2.31335 net_r[141] <= net_w[141];
end
always @(posedge net_w[142] or negedge net_w[142]) begin
	#1.47213 net_r[142] <= net_w[142];
end
always @(posedge net_w[143] or negedge net_w[143]) begin
	#2.31335 net_r[143] <= net_w[143];
end
always @(posedge net_w[144] or negedge net_w[144]) begin
	#1.68244 net_r[144] <= net_w[144];
end
always @(posedge net_w[145] or negedge net_w[145]) begin
	#1.89274 net_r[145] <= net_w[145];
end
always @(posedge net_w[146] or negedge net_w[146]) begin
	#1.05152 net_r[146] <= net_w[146];
end
always @(posedge net_w[147] or negedge net_w[147]) begin
	#1.78759 net_r[147] <= net_w[147];
end
always @(posedge net_w[148] or negedge net_w[148]) begin
	#1.57729 net_r[148] <= net_w[148];
end
always @(posedge net_w[149] or negedge net_w[149]) begin
	#2.52366 net_r[149] <= net_w[149];
end
always @(posedge net_w[150] or negedge net_w[150]) begin
	#1.47213 net_r[150] <= net_w[150];
end
always @(posedge net_w[151] or negedge net_w[151]) begin
	#2.10305 net_r[151] <= net_w[151];
end
always @(posedge net_w[152] or negedge net_w[152]) begin
	#1.47213 net_r[152] <= net_w[152];
end
always @(posedge net_w[153] or negedge net_w[153]) begin
	#2.31335 net_r[153] <= net_w[153];
end
always @(posedge net_w[154] or negedge net_w[154]) begin
	#1.36698 net_r[154] <= net_w[154];
end
always @(posedge net_w[155] or negedge net_w[155]) begin
	#2.31335 net_r[155] <= net_w[155];
end
always @(posedge net_w[156] or negedge net_w[156]) begin
	#1.57729 net_r[156] <= net_w[156];
end
always @(posedge net_w[157] or negedge net_w[157]) begin
	#1.9979 net_r[157] <= net_w[157];
end
always @(posedge net_w[158] or negedge net_w[158]) begin
	#0.946372 net_r[158] <= net_w[158];
end
always @(posedge net_w[159] or negedge net_w[159]) begin
	#1.9979 net_r[159] <= net_w[159];
end
always @(posedge net_w[160] or negedge net_w[160]) begin
	#1.57729 net_r[160] <= net_w[160];
end
always @(posedge net_w[161] or negedge net_w[161]) begin
	#2.41851 net_r[161] <= net_w[161];
end
always @(posedge net_w[162] or negedge net_w[162]) begin
	#1.26183 net_r[162] <= net_w[162];
end
always @(posedge net_w[163] or negedge net_w[163]) begin
	#2.52366 net_r[163] <= net_w[163];
end
always @(posedge net_w[164] or negedge net_w[164]) begin
	#1.47213 net_r[164] <= net_w[164];
end
always @(posedge net_w[165] or negedge net_w[165]) begin
	#2.10305 net_r[165] <= net_w[165];
end
always @(posedge net_w[166] or negedge net_w[166]) begin
	#1.47213 net_r[166] <= net_w[166];
end
always @(posedge net_w[167] or negedge net_w[167]) begin
	#2.2082 net_r[167] <= net_w[167];
end
always @(posedge net_w[168] or negedge net_w[168]) begin
	#1.36698 net_r[168] <= net_w[168];
end
always @(posedge net_w[169] or negedge net_w[169]) begin
	#2.31335 net_r[169] <= net_w[169];
end
always @(posedge net_w[170] or negedge net_w[170]) begin
	#1.47213 net_r[170] <= net_w[170];
end
always @(posedge net_w[171] or negedge net_w[171]) begin
	#2.10305 net_r[171] <= net_w[171];
end
always @(posedge net_w[172] or negedge net_w[172]) begin
	#1.05152 net_r[172] <= net_w[172];
end
always @(posedge net_w[173] or negedge net_w[173]) begin
	#1.78759 net_r[173] <= net_w[173];
end
always @(posedge net_w[174] or negedge net_w[174]) begin
	#1.47213 net_r[174] <= net_w[174];
end
always @(posedge net_w[175] or negedge net_w[175]) begin
	#1.36698 net_r[175] <= net_w[175];
end
always @(posedge net_w[176] or negedge net_w[176]) begin
	#1.26183 net_r[176] <= net_w[176];
end
always @(posedge net_w[177] or negedge net_w[177]) begin
	#2.31335 net_r[177] <= net_w[177];
end
always @(posedge net_w[178] or negedge net_w[178]) begin
	#0.946372 net_r[178] <= net_w[178];
end
always @(posedge net_w[179] or negedge net_w[179]) begin
	#3.47003 net_r[179] <= net_w[179];
end
always @(posedge net_w[180] or negedge net_w[180]) begin
	#7.04522 net_r[180] <= net_w[180];
end
always @(posedge net_w[181] or negedge net_w[181]) begin
	#5.36278 net_r[181] <= net_w[181];
end
always @(posedge net_w[182] or negedge net_w[182]) begin
	#4.10095 net_r[182] <= net_w[182];
end
always @(posedge net_w[183] or negedge net_w[183]) begin
	#2.52366 net_r[183] <= net_w[183];
end
always @(posedge net_w[184] or negedge net_w[184]) begin
	#2.94427 net_r[184] <= net_w[184];
end
always @(posedge net_w[185] or negedge net_w[185]) begin
	#3.15457 net_r[185] <= net_w[185];
end
always @(posedge net_w[186] or negedge net_w[186]) begin
	#2.2082 net_r[186] <= net_w[186];
end
always @(posedge net_w[187] or negedge net_w[187]) begin
	#2.41851 net_r[187] <= net_w[187];
end
always @(posedge net_w[188] or negedge net_w[188]) begin
	#1.57729 net_r[188] <= net_w[188];
end
always @(posedge net_w[189] or negedge net_w[189]) begin
	#2.94427 net_r[189] <= net_w[189];
end
always @(posedge net_w[190] or negedge net_w[190]) begin
	#1.15668 net_r[190] <= net_w[190];
end
always @(posedge net_w[191] or negedge net_w[191]) begin
	#2.10305 net_r[191] <= net_w[191];
end
always @(posedge net_w[192] or negedge net_w[192]) begin
	#1.26183 net_r[192] <= net_w[192];
end
always @(posedge net_w[193] or negedge net_w[193]) begin
	#2.31335 net_r[193] <= net_w[193];
end
always @(posedge net_w[194] or negedge net_w[194]) begin
	#1.26183 net_r[194] <= net_w[194];
end
always @(posedge net_w[195] or negedge net_w[195]) begin
	#2.41851 net_r[195] <= net_w[195];
end
always @(posedge net_w[196] or negedge net_w[196]) begin
	#2.10305 net_r[196] <= net_w[196];
end
always @(posedge net_w[197] or negedge net_w[197]) begin
	#1.89274 net_r[197] <= net_w[197];
end
always @(posedge net_w[198] or negedge net_w[198]) begin
	#1.9979 net_r[198] <= net_w[198];
end
always @(posedge net_w[199] or negedge net_w[199]) begin
	#2.31335 net_r[199] <= net_w[199];
end
always @(posedge net_w[200] or negedge net_w[200]) begin
	#2.83912 net_r[200] <= net_w[200];
end
always @(posedge net_w[201] or negedge net_w[201]) begin
	#3.47003 net_r[201] <= net_w[201];
end
always @(posedge net_w[202] or negedge net_w[202]) begin
	#1.9979 net_r[202] <= net_w[202];
end
always @(posedge net_w[203] or negedge net_w[203]) begin
	#2.41851 net_r[203] <= net_w[203];
end
always @(posedge net_w[204] or negedge net_w[204]) begin
	#1.68244 net_r[204] <= net_w[204];
end
always @(posedge net_w[205] or negedge net_w[205]) begin
	#2.73396 net_r[205] <= net_w[205];
end
always @(posedge net_w[206] or negedge net_w[206]) begin
	#0.946372 net_r[206] <= net_w[206];
end
always @(posedge net_w[207] or negedge net_w[207]) begin
	#1.9979 net_r[207] <= net_w[207];
end
always @(posedge net_w[208] or negedge net_w[208]) begin
	#1.15668 net_r[208] <= net_w[208];
end
always @(posedge net_w[209] or negedge net_w[209]) begin
	#2.31335 net_r[209] <= net_w[209];
end
always @(posedge net_w[210] or negedge net_w[210]) begin
	#1.26183 net_r[210] <= net_w[210];
end
always @(posedge net_w[211] or negedge net_w[211]) begin
	#2.41851 net_r[211] <= net_w[211];
end
always @(posedge net_w[212] or negedge net_w[212]) begin
	#4.62671 net_r[212] <= net_w[212];
end
always @(posedge net_w[213] or negedge net_w[213]) begin
	#2.31335 net_r[213] <= net_w[213];
end
always @(posedge net_w[214] or negedge net_w[214]) begin
	#2.73396 net_r[214] <= net_w[214];
end
always @(posedge net_w[215] or negedge net_w[215]) begin
	#3.89064 net_r[215] <= net_w[215];
end
always @(posedge net_w[216] or negedge net_w[216]) begin
	#1.78759 net_r[216] <= net_w[216];
end
always @(posedge net_w[217] or negedge net_w[217]) begin
	#2.52366 net_r[217] <= net_w[217];
end
always @(posedge net_w[218] or negedge net_w[218]) begin
	#1.78759 net_r[218] <= net_w[218];
end
always @(posedge net_w[219] or negedge net_w[219]) begin
	#2.62881 net_r[219] <= net_w[219];
end
always @(posedge net_w[220] or negedge net_w[220]) begin
	#1.05152 net_r[220] <= net_w[220];
end
always @(posedge net_w[221] or negedge net_w[221]) begin
	#1.9979 net_r[221] <= net_w[221];
end
always @(posedge net_w[222] or negedge net_w[222]) begin
	#1.36698 net_r[222] <= net_w[222];
end
always @(posedge net_w[223] or negedge net_w[223]) begin
	#5.46793 net_r[223] <= net_w[223];
end
always @(posedge net_w[224] or negedge net_w[224]) begin
	#3.89064 net_r[224] <= net_w[224];
end
always @(posedge net_w[225] or negedge net_w[225]) begin
	#2.2082 net_r[225] <= net_w[225];
end
always @(posedge net_w[226] or negedge net_w[226]) begin
	#2.52366 net_r[226] <= net_w[226];
end
always @(posedge net_w[227] or negedge net_w[227]) begin
	#4.10095 net_r[227] <= net_w[227];
end
always @(posedge net_w[228] or negedge net_w[228]) begin
	#1.47213 net_r[228] <= net_w[228];
end
always @(posedge net_w[229] or negedge net_w[229]) begin
	#2.62881 net_r[229] <= net_w[229];
end
always @(posedge net_w[230] or negedge net_w[230]) begin
	#1.78759 net_r[230] <= net_w[230];
end
always @(posedge net_w[231] or negedge net_w[231]) begin
	#2.52366 net_r[231] <= net_w[231];
end
always @(posedge net_w[232] or negedge net_w[232]) begin
	#3.57518 net_r[232] <= net_w[232];
end
always @(posedge net_w[233] or negedge net_w[233]) begin
	#5.25762 net_r[233] <= net_w[233];
end
always @(posedge net_w[234] or negedge net_w[234]) begin
	#3.15457 net_r[234] <= net_w[234];
end
always @(posedge net_w[235] or negedge net_w[235]) begin
	#2.2082 net_r[235] <= net_w[235];
end
always @(posedge net_w[236] or negedge net_w[236]) begin
	#2.41851 net_r[236] <= net_w[236];
end
always @(posedge net_w[237] or negedge net_w[237]) begin
	#4.52156 net_r[237] <= net_w[237];
end
always @(posedge net_w[238] or negedge net_w[238]) begin
	#1.57729 net_r[238] <= net_w[238];
end
always @(posedge net_w[239] or negedge net_w[239]) begin
	#4.62671 net_r[239] <= net_w[239];
end
always @(posedge net_w[240] or negedge net_w[240]) begin
	#2.94427 net_r[240] <= net_w[240];
end
always @(posedge net_w[241] or negedge net_w[241]) begin
	#5.46793 net_r[241] <= net_w[241];
end
always @(posedge net_w[242] or negedge net_w[242]) begin
	#2.41851 net_r[242] <= net_w[242];
end
always @(posedge net_w[243] or negedge net_w[243]) begin
	#2.31335 net_r[243] <= net_w[243];
end
always @(posedge net_w[244] or negedge net_w[244]) begin
	#3.68034 net_r[244] <= net_w[244];
end
always @(posedge net_w[245] or negedge net_w[245]) begin
	#3.78549 net_r[245] <= net_w[245];
end
always @(posedge net_w[246] or negedge net_w[246]) begin
	#2.62881 net_r[246] <= net_w[246];
end
always @(posedge net_w[247] or negedge net_w[247]) begin
	#6.72976 net_r[247] <= net_w[247];
end
always @(posedge net_w[248] or negedge net_w[248]) begin
	#1.89274 net_r[248] <= net_w[248];
end
always @(posedge net_w[249] or negedge net_w[249]) begin
	#2.2082 net_r[249] <= net_w[249];
end
always @(posedge net_w[250] or negedge net_w[250]) begin
	#1.68244 net_r[250] <= net_w[250];
end
always @(posedge net_w[251] or negedge net_w[251]) begin
	#2.94427 net_r[251] <= net_w[251];
end
always @(posedge net_w[252] or negedge net_w[252]) begin
	#2.73396 net_r[252] <= net_w[252];
end
always @(posedge net_w[253] or negedge net_w[253]) begin
	#2.31335 net_r[253] <= net_w[253];
end
always @(posedge net_w[254] or negedge net_w[254]) begin
	#3.25973 net_r[254] <= net_w[254];
end
always @(posedge net_w[255] or negedge net_w[255]) begin
	#2.62881 net_r[255] <= net_w[255];
end
always @(posedge net_w[256] or negedge net_w[256]) begin
	#0.84122 net_r[256] <= net_w[256];
end
always @(posedge net_w[257] or negedge net_w[257]) begin
	#2.31335 net_r[257] <= net_w[257];
end
always @(posedge net_w[258] or negedge net_w[258]) begin
	#1.57729 net_r[258] <= net_w[258];
end
always @(posedge net_w[259] or negedge net_w[259]) begin
	#2.52366 net_r[259] <= net_w[259];
end
always @(posedge net_w[260] or negedge net_w[260]) begin
	#1.9979 net_r[260] <= net_w[260];
end
always @(posedge net_w[261] or negedge net_w[261]) begin
	#1.78759 net_r[261] <= net_w[261];
end
always @(posedge net_w[262] or negedge net_w[262]) begin
	#1.9979 net_r[262] <= net_w[262];
end
always @(posedge net_w[263] or negedge net_w[263]) begin
	#1.15668 net_r[263] <= net_w[263];
end
always @(posedge net_w[264] or negedge net_w[264]) begin
	#4.31125 net_r[264] <= net_w[264];
end
always @(posedge net_w[265] or negedge net_w[265]) begin
	#3.57518 net_r[265] <= net_w[265];
end
always @(posedge net_w[266] or negedge net_w[266]) begin
	#1.26183 net_r[266] <= net_w[266];
end
always @(posedge net_w[267] or negedge net_w[267]) begin
	#3.68034 net_r[267] <= net_w[267];
end
always @(posedge net_w[268] or negedge net_w[268]) begin
	#2.94427 net_r[268] <= net_w[268];
end
always @(posedge net_w[269] or negedge net_w[269]) begin
	#4.10095 net_r[269] <= net_w[269];
end
always @(posedge net_w[270] or negedge net_w[270]) begin
	#3.25973 net_r[270] <= net_w[270];
end
always @(posedge net_w[271] or negedge net_w[271]) begin
	#0.736067 net_r[271] <= net_w[271];
end
always @(posedge net_w[272] or negedge net_w[272]) begin
	#2.83912 net_r[272] <= net_w[272];
end
always @(posedge net_w[273] or negedge net_w[273]) begin
	#1.9979 net_r[273] <= net_w[273];
end
always @(posedge net_w[274] or negedge net_w[274]) begin
	#3.25973 net_r[274] <= net_w[274];
end
always @(posedge net_w[275] or negedge net_w[275]) begin
	#2.41851 net_r[275] <= net_w[275];
end
always @(posedge net_w[276] or negedge net_w[276]) begin
	#1.57729 net_r[276] <= net_w[276];
end
always @(posedge net_w[277] or negedge net_w[277]) begin
	#2.31335 net_r[277] <= net_w[277];
end
always @(posedge net_w[278] or negedge net_w[278]) begin
	#1.36698 net_r[278] <= net_w[278];
end
always @(posedge net_w[279] or negedge net_w[279]) begin
	#9.77918 net_r[279] <= net_w[279];
end
always @(posedge net_w[280] or negedge net_w[280]) begin
	#7.46583 net_r[280] <= net_w[280];
end
always @(posedge net_w[281] or negedge net_w[281]) begin
	#8.30705 net_r[281] <= net_w[281];
end
always @(posedge net_w[282] or negedge net_w[282]) begin
	#7.36067 net_r[282] <= net_w[282];
end
always @(posedge net_w[283] or negedge net_w[283]) begin
	#9.98948 net_r[283] <= net_w[283];
end
always @(posedge net_w[284] or negedge net_w[284]) begin
	#7.57098 net_r[284] <= net_w[284];
end
always @(posedge net_w[285] or negedge net_w[285]) begin
	#2.2082 net_r[285] <= net_w[285];
end
always @(posedge net_w[286] or negedge net_w[286]) begin
	#1.68244 net_r[286] <= net_w[286];
end
always @(posedge net_w[287] or negedge net_w[287]) begin
	#8.09674 net_r[287] <= net_w[287];
end
always @(posedge net_w[288] or negedge net_w[288]) begin
	#4.31125 net_r[288] <= net_w[288];
end
always @(posedge net_w[289] or negedge net_w[289]) begin
	#6.09884 net_r[289] <= net_w[289];
end
always @(posedge net_w[290] or negedge net_w[290]) begin
	#1.89274 net_r[290] <= net_w[290];
end
always @(posedge net_w[291] or negedge net_w[291]) begin
	#1.26183 net_r[291] <= net_w[291];
end
always @(posedge net_w[292] or negedge net_w[292]) begin
	#7.57098 net_r[292] <= net_w[292];
end
always @(posedge net_w[293] or negedge net_w[293]) begin
	#3.57518 net_r[293] <= net_w[293];
end
always @(posedge net_w[294] or negedge net_w[294]) begin
	#5.67823 net_r[294] <= net_w[294];
end
always @(posedge net_w[295] or negedge net_w[295]) begin
	#2.62881 net_r[295] <= net_w[295];
end
always @(posedge net_w[296] or negedge net_w[296]) begin
	#1.89274 net_r[296] <= net_w[296];
end
always @(posedge net_w[297] or negedge net_w[297]) begin
	#4.94217 net_r[297] <= net_w[297];
end
always @(posedge net_w[298] or negedge net_w[298]) begin
	#1.57729 net_r[298] <= net_w[298];
end
always @(posedge net_w[299] or negedge net_w[299]) begin
	#3.25973 net_r[299] <= net_w[299];
end
always @(posedge net_w[300] or negedge net_w[300]) begin
	#2.62881 net_r[300] <= net_w[300];
end
always @(posedge net_w[301] or negedge net_w[301]) begin
	#1.78759 net_r[301] <= net_w[301];
end
always @(posedge net_w[302] or negedge net_w[302]) begin
	#4.94217 net_r[302] <= net_w[302];
end
always @(posedge net_w[303] or negedge net_w[303]) begin
	#1.26183 net_r[303] <= net_w[303];
end
always @(posedge net_w[304] or negedge net_w[304]) begin
	#2.83912 net_r[304] <= net_w[304];
end
always @(posedge net_w[305] or negedge net_w[305]) begin
	#2.2082 net_r[305] <= net_w[305];
end
always @(posedge net_w[306] or negedge net_w[306]) begin
	#1.36698 net_r[306] <= net_w[306];
end
always @(posedge net_w[307] or negedge net_w[307]) begin
	#4.62671 net_r[307] <= net_w[307];
end
always @(posedge net_w[308] or negedge net_w[308]) begin
	#0.42061 net_r[308] <= net_w[308];
end
always @(posedge net_w[309] or negedge net_w[309]) begin
	#2.10305 net_r[309] <= net_w[309];
end
always @(posedge net_w[310] or negedge net_w[310]) begin
	#17.3502 net_r[310] <= net_w[310];
end
always @(posedge net_w[311] or negedge net_w[311]) begin
	#16.6141 net_r[311] <= net_w[311];
end
always @(posedge net_w[312] or negedge net_w[312]) begin
	#1.89274 net_r[312] <= net_w[312];
end
always @(posedge net_w[313] or negedge net_w[313]) begin
	#2.73396 net_r[313] <= net_w[313];
end
always @(posedge net_w[314] or negedge net_w[314]) begin
	#1.05152 net_r[314] <= net_w[314];
end
always @(posedge net_w[315] or negedge net_w[315]) begin
	#1.26183 net_r[315] <= net_w[315];
end
always @(posedge net_w[316] or negedge net_w[316]) begin
	#4.10095 net_r[316] <= net_w[316];
end
always @(posedge net_w[317] or negedge net_w[317]) begin
	#2.94427 net_r[317] <= net_w[317];
end
always @(posedge net_w[318] or negedge net_w[318]) begin
	#5.67823 net_r[318] <= net_w[318];
end
always @(posedge net_w[319] or negedge net_w[319]) begin
	#4.83701 net_r[319] <= net_w[319];
end
always @(posedge net_w[320] or negedge net_w[320]) begin
	#1.78759 net_r[320] <= net_w[320];
end
always @(posedge net_w[321] or negedge net_w[321]) begin
	#2.94427 net_r[321] <= net_w[321];
end
always @(posedge net_w[322] or negedge net_w[322]) begin
	#1.26183 net_r[322] <= net_w[322];
end
always @(posedge net_w[323] or negedge net_w[323]) begin
	#3.89064 net_r[323] <= net_w[323];
end
always @(posedge net_w[324] or negedge net_w[324]) begin
	#2.10305 net_r[324] <= net_w[324];
end
always @(posedge net_w[325] or negedge net_w[325]) begin
	#2.94427 net_r[325] <= net_w[325];
end
always @(posedge net_w[326] or negedge net_w[326]) begin
	#1.78759 net_r[326] <= net_w[326];
end
always @(posedge net_w[327] or negedge net_w[327]) begin
	#2.31335 net_r[327] <= net_w[327];
end
always @(posedge net_w[328] or negedge net_w[328]) begin
	#5.04732 net_r[328] <= net_w[328];
end
always @(posedge net_w[329] or negedge net_w[329]) begin
	#1.36698 net_r[329] <= net_w[329];
end
always @(posedge net_w[330] or negedge net_w[330]) begin
	#3.99579 net_r[330] <= net_w[330];
end
always @(posedge net_w[331] or negedge net_w[331]) begin
	#1.36698 net_r[331] <= net_w[331];
end
always @(posedge net_w[332] or negedge net_w[332]) begin
	#17.4553 net_r[332] <= net_w[332];
end
always @(posedge net_w[333] or negedge net_w[333]) begin
	#1.26183 net_r[333] <= net_w[333];
end
always @(posedge net_w[334] or negedge net_w[334]) begin
	#2.83912 net_r[334] <= net_w[334];
end
always @(posedge net_w[335] or negedge net_w[335]) begin
	#0.630915 net_r[335] <= net_w[335];
end
always @(posedge net_w[336] or negedge net_w[336]) begin
	#2.31335 net_r[336] <= net_w[336];
end
always @(posedge net_w[337] or negedge net_w[337]) begin
	#0.736067 net_r[337] <= net_w[337];
end
always @(posedge net_w[338] or negedge net_w[338]) begin
	#2.41851 net_r[338] <= net_w[338];
end
always @(posedge net_w[339] or negedge net_w[339]) begin
	#0.630915 net_r[339] <= net_w[339];
end
always @(posedge net_w[340] or negedge net_w[340]) begin
	#2.10305 net_r[340] <= net_w[340];
end
always @(posedge net_w[341] or negedge net_w[341]) begin
	#0.525762 net_r[341] <= net_w[341];
end
always @(posedge net_w[342] or negedge net_w[342]) begin
	#1.9979 net_r[342] <= net_w[342];
end
always @(posedge net_w[343] or negedge net_w[343]) begin
	#0.42061 net_r[343] <= net_w[343];
end
always @(posedge net_w[344] or negedge net_w[344]) begin
	#1.89274 net_r[344] <= net_w[344];
end
always @(posedge net_w[345] or negedge net_w[345]) begin
	#0.525762 net_r[345] <= net_w[345];
end
always @(posedge net_w[346] or negedge net_w[346]) begin
	#1.78759 net_r[346] <= net_w[346];
end
always @(posedge net_w[347] or negedge net_w[347]) begin
	#0.630915 net_r[347] <= net_w[347];
end
always @(posedge net_w[348] or negedge net_w[348]) begin
	#0.946372 net_r[348] <= net_w[348];
end
always @(posedge net_w[349] or negedge net_w[349]) begin
	#1.47213 net_r[349] <= net_w[349];
end
always @(posedge net_w[350] or negedge net_w[350]) begin
	#0.84122 net_r[350] <= net_w[350];
end
always @(posedge net_w[351] or negedge net_w[351]) begin
	#1.57729 net_r[351] <= net_w[351];
end
always @(posedge net_w[352] or negedge net_w[352]) begin
	#0.736067 net_r[352] <= net_w[352];
end
always @(posedge net_w[353] or negedge net_w[353]) begin
	#1.47213 net_r[353] <= net_w[353];
end
always @(posedge net_w[354] or negedge net_w[354]) begin
	#0.630915 net_r[354] <= net_w[354];
end
always @(posedge net_w[355] or negedge net_w[355]) begin
	#1.57729 net_r[355] <= net_w[355];
end
always @(posedge net_w[356] or negedge net_w[356]) begin
	#0.525762 net_r[356] <= net_w[356];
end
always @(posedge net_w[357] or negedge net_w[357]) begin
	#1.47213 net_r[357] <= net_w[357];
end
always @(posedge net_w[358] or negedge net_w[358]) begin
	#0.42061 net_r[358] <= net_w[358];
end
always @(posedge net_w[359] or negedge net_w[359]) begin
	#1.57729 net_r[359] <= net_w[359];
end
always @(posedge net_w[360] or negedge net_w[360]) begin
	#0.525762 net_r[360] <= net_w[360];
end
always @(posedge net_w[361] or negedge net_w[361]) begin
	#1.68244 net_r[361] <= net_w[361];
end
always @(posedge net_w[362] or negedge net_w[362]) begin
	#0.630915 net_r[362] <= net_w[362];
end
always @(posedge net_w[363] or negedge net_w[363]) begin
	#1.78759 net_r[363] <= net_w[363];
end
always @(posedge net_w[364] or negedge net_w[364]) begin
	#1.9979 net_r[364] <= net_w[364];
end
always @(posedge net_w[365] or negedge net_w[365]) begin
	#2.62881 net_r[365] <= net_w[365];
end
always @(posedge net_w[366] or negedge net_w[366]) begin
	#1.36698 net_r[366] <= net_w[366];
end
always @(posedge net_w[367] or negedge net_w[367]) begin
	#2.83912 net_r[367] <= net_w[367];
end
always @(posedge net_w[368] or negedge net_w[368]) begin
	#2.41851 net_r[368] <= net_w[368];
end
always @(posedge net_w[369] or negedge net_w[369]) begin
	#2.31335 net_r[369] <= net_w[369];
end
always @(posedge net_w[370] or negedge net_w[370]) begin
	#2.31335 net_r[370] <= net_w[370];
end
always @(posedge net_w[371] or negedge net_w[371]) begin
	#2.10305 net_r[371] <= net_w[371];
end
always @(posedge net_w[372] or negedge net_w[372]) begin
	#2.31335 net_r[372] <= net_w[372];
end
always @(posedge net_w[373] or negedge net_w[373]) begin
	#2.2082 net_r[373] <= net_w[373];
end
always @(posedge net_w[374] or negedge net_w[374]) begin
	#2.41851 net_r[374] <= net_w[374];
end
always @(posedge net_w[375] or negedge net_w[375]) begin
	#1.89274 net_r[375] <= net_w[375];
end
always @(posedge net_w[376] or negedge net_w[376]) begin
	#2.10305 net_r[376] <= net_w[376];
end
always @(posedge net_w[377] or negedge net_w[377]) begin
	#1.57729 net_r[377] <= net_w[377];
end
always @(posedge net_w[378] or negedge net_w[378]) begin
	#1.57729 net_r[378] <= net_w[378];
end
always @(posedge net_w[379] or negedge net_w[379]) begin
	#0.946372 net_r[379] <= net_w[379];
end
always @(posedge net_w[380] or negedge net_w[380]) begin
	#0.946372 net_r[380] <= net_w[380];
end
always @(posedge net_w[381] or negedge net_w[381]) begin
	#1.68244 net_r[381] <= net_w[381];
end
always @(posedge net_w[382] or negedge net_w[382]) begin
	#0.525762 net_r[382] <= net_w[382];
end
always @(posedge net_w[383] or negedge net_w[383]) begin
	#1.36698 net_r[383] <= net_w[383];
end
always @(posedge net_w[384] or negedge net_w[384]) begin
	#1.15668 net_r[384] <= net_w[384];
end
always @(posedge net_w[385] or negedge net_w[385]) begin
	#1.68244 net_r[385] <= net_w[385];
end
always @(posedge net_w[386] or negedge net_w[386]) begin
	#1.47213 net_r[386] <= net_w[386];
end
always @(posedge net_w[387] or negedge net_w[387]) begin
	#1.89274 net_r[387] <= net_w[387];
end
always @(posedge net_w[388] or negedge net_w[388]) begin
	#1.57729 net_r[388] <= net_w[388];
end
always @(posedge net_w[389] or negedge net_w[389]) begin
	#1.89274 net_r[389] <= net_w[389];
end
always @(posedge net_w[390] or negedge net_w[390]) begin
	#1.15668 net_r[390] <= net_w[390];
end
always @(posedge net_w[391] or negedge net_w[391]) begin
	#1.36698 net_r[391] <= net_w[391];
end
always @(posedge net_w[392] or negedge net_w[392]) begin
	#0.736067 net_r[392] <= net_w[392];
end
always @(posedge net_w[393] or negedge net_w[393]) begin
	#1.47213 net_r[393] <= net_w[393];
end
always @(posedge net_w[394] or negedge net_w[394]) begin
	#1.15668 net_r[394] <= net_w[394];
end
always @(posedge net_w[395] or negedge net_w[395]) begin
	#1.9979 net_r[395] <= net_w[395];
end
always @(posedge net_w[396] or negedge net_w[396]) begin
	#2.52366 net_r[396] <= net_w[396];
end
always @(posedge net_w[397] or negedge net_w[397]) begin
	#2.10305 net_r[397] <= net_w[397];
end
always @(posedge net_w[398] or negedge net_w[398]) begin
	#1.89274 net_r[398] <= net_w[398];
end
always @(posedge net_w[399] or negedge net_w[399]) begin
	#2.2082 net_r[399] <= net_w[399];
end
always @(posedge net_w[400] or negedge net_w[400]) begin
	#2.52366 net_r[400] <= net_w[400];
end
always @(posedge net_w[401] or negedge net_w[401]) begin
	#2.52366 net_r[401] <= net_w[401];
end
always @(posedge net_w[402] or negedge net_w[402]) begin
	#2.52366 net_r[402] <= net_w[402];
end
always @(posedge net_w[403] or negedge net_w[403]) begin
	#1.9979 net_r[403] <= net_w[403];
end
always @(posedge net_w[404] or negedge net_w[404]) begin
	#2.83912 net_r[404] <= net_w[404];
end
always @(posedge net_w[405] or negedge net_w[405]) begin
	#0.630915 net_r[405] <= net_w[405];
end
always @(posedge net_w[406] or negedge net_w[406]) begin
	#1.89274 net_r[406] <= net_w[406];
end
always @(posedge net_w[407] or negedge net_w[407]) begin
	#2.10305 net_r[407] <= net_w[407];
end
always @(posedge net_w[408] or negedge net_w[408]) begin
	#3.68034 net_r[408] <= net_w[408];
end
always @(posedge net_w[409] or negedge net_w[409]) begin
	#2.2082 net_r[409] <= net_w[409];
end
always @(posedge net_w[410] or negedge net_w[410]) begin
	#1.36698 net_r[410] <= net_w[410];
end
always @(posedge net_w[411] or negedge net_w[411]) begin
	#3.47003 net_r[411] <= net_w[411];
end
always @(posedge net_w[412] or negedge net_w[412]) begin
	#0.84122 net_r[412] <= net_w[412];
end
always @(posedge net_w[413] or negedge net_w[413]) begin
	#3.78549 net_r[413] <= net_w[413];
end
always @(posedge net_w[414] or negedge net_w[414]) begin
	#0.946372 net_r[414] <= net_w[414];
end
always @(posedge net_w[415] or negedge net_w[415]) begin
	#3.15457 net_r[415] <= net_w[415];
end
always @(posedge net_w[416] or negedge net_w[416]) begin
	#0.525762 net_r[416] <= net_w[416];
end
always @(posedge net_w[417] or negedge net_w[417]) begin
	#2.73396 net_r[417] <= net_w[417];
end
always @(posedge net_w[418] or negedge net_w[418]) begin
	#1.89274 net_r[418] <= net_w[418];
end
always @(posedge net_w[419] or negedge net_w[419]) begin
	#1.78759 net_r[419] <= net_w[419];
end
always @(posedge net_w[420] or negedge net_w[420]) begin
	#1.15668 net_r[420] <= net_w[420];
end
always @(posedge net_w[421] or negedge net_w[421]) begin
	#1.57729 net_r[421] <= net_w[421];
end
always @(posedge net_w[422] or negedge net_w[422]) begin
	#1.26183 net_r[422] <= net_w[422];
end
always @(posedge net_w[423] or negedge net_w[423]) begin
	#1.89274 net_r[423] <= net_w[423];
end
always @(posedge net_w[424] or negedge net_w[424]) begin
	#0.630915 net_r[424] <= net_w[424];
end
always @(posedge net_w[425] or negedge net_w[425]) begin
	#1.57729 net_r[425] <= net_w[425];
end
always @(posedge net_w[426] or negedge net_w[426]) begin
	#1.05152 net_r[426] <= net_w[426];
end
always @(posedge net_w[427] or negedge net_w[427]) begin
	#1.9979 net_r[427] <= net_w[427];
end
always @(posedge net_w[428] or negedge net_w[428]) begin
	#0.946372 net_r[428] <= net_w[428];
end
always @(posedge net_w[429] or negedge net_w[429]) begin
	#1.9979 net_r[429] <= net_w[429];
end
always @(posedge net_w[430] or negedge net_w[430]) begin
	#1.36698 net_r[430] <= net_w[430];
end
always @(posedge net_w[431] or negedge net_w[431]) begin
	#2.2082 net_r[431] <= net_w[431];
end
always @(posedge net_w[432] or negedge net_w[432]) begin
	#1.47213 net_r[432] <= net_w[432];
end
always @(posedge net_w[433] or negedge net_w[433]) begin
	#2.31335 net_r[433] <= net_w[433];
end
always @(posedge net_w[434] or negedge net_w[434]) begin
	#1.89274 net_r[434] <= net_w[434];
end
always @(posedge net_w[435] or negedge net_w[435]) begin
	#0.42061 net_r[435] <= net_w[435];
end
always @(posedge net_w[436] or negedge net_w[436]) begin
	#2.31335 net_r[436] <= net_w[436];
end
always @(posedge net_w[437] or negedge net_w[437]) begin
	#0.630915 net_r[437] <= net_w[437];
end
always @(posedge net_w[438] or negedge net_w[438]) begin
	#2.10305 net_r[438] <= net_w[438];
end
always @(posedge net_w[439] or negedge net_w[439]) begin
	#0.736067 net_r[439] <= net_w[439];
end
always @(posedge net_w[440] or negedge net_w[440]) begin
	#1.89274 net_r[440] <= net_w[440];
end
always @(posedge net_w[441] or negedge net_w[441]) begin
	#0.84122 net_r[441] <= net_w[441];
end
always @(posedge net_w[442] or negedge net_w[442]) begin
	#1.89274 net_r[442] <= net_w[442];
end
always @(posedge net_w[443] or negedge net_w[443]) begin
	#1.15668 net_r[443] <= net_w[443];
end
always @(posedge net_w[444] or negedge net_w[444]) begin
	#2.10305 net_r[444] <= net_w[444];
end
always @(posedge net_w[445] or negedge net_w[445]) begin
	#1.36698 net_r[445] <= net_w[445];
end
always @(posedge net_w[446] or negedge net_w[446]) begin
	#0.630915 net_r[446] <= net_w[446];
end
always @(posedge net_w[447] or negedge net_w[447]) begin
	#1.78759 net_r[447] <= net_w[447];
end
always @(posedge net_w[448] or negedge net_w[448]) begin
	#1.68244 net_r[448] <= net_w[448];
end
always @(posedge net_w[449] or negedge net_w[449]) begin
	#1.78759 net_r[449] <= net_w[449];
end
always @(posedge net_w[450] or negedge net_w[450]) begin
	#1.47213 net_r[450] <= net_w[450];
end
always @(posedge net_w[451] or negedge net_w[451]) begin
	#1.47213 net_r[451] <= net_w[451];
end
always @(posedge net_w[452] or negedge net_w[452]) begin
	#1.68244 net_r[452] <= net_w[452];
end
always @(posedge net_w[453] or negedge net_w[453]) begin
	#1.57729 net_r[453] <= net_w[453];
end
always @(posedge net_w[454] or negedge net_w[454]) begin
	#3.25973 net_r[454] <= net_w[454];
end
always @(posedge net_w[455] or negedge net_w[455]) begin
	#3.15457 net_r[455] <= net_w[455];
end
always @(posedge net_w[456] or negedge net_w[456]) begin
	#3.47003 net_r[456] <= net_w[456];
end
always @(posedge net_w[457] or negedge net_w[457]) begin
	#3.47003 net_r[457] <= net_w[457];
end
always @(posedge net_w[458] or negedge net_w[458]) begin
	#2.73396 net_r[458] <= net_w[458];
end
always @(posedge net_w[459] or negedge net_w[459]) begin
	#1.78759 net_r[459] <= net_w[459];
end
always @(posedge net_w[460] or negedge net_w[460]) begin
	#2.52366 net_r[460] <= net_w[460];
end
always @(posedge net_w[461] or negedge net_w[461]) begin
	#1.36698 net_r[461] <= net_w[461];
end
always @(posedge net_w[462] or negedge net_w[462]) begin
	#1.9979 net_r[462] <= net_w[462];
end
always @(posedge net_w[463] or negedge net_w[463]) begin
	#1.26183 net_r[463] <= net_w[463];
end
always @(posedge net_w[464] or negedge net_w[464]) begin
	#1.78759 net_r[464] <= net_w[464];
end
always @(posedge net_w[465] or negedge net_w[465]) begin
	#1.05152 net_r[465] <= net_w[465];
end
always @(posedge net_w[466] or negedge net_w[466]) begin
	#1.9979 net_r[466] <= net_w[466];
end
always @(posedge net_w[467] or negedge net_w[467]) begin
	#1.15668 net_r[467] <= net_w[467];
end
always @(posedge net_w[468] or negedge net_w[468]) begin
	#2.31335 net_r[468] <= net_w[468];
end
always @(posedge net_w[469] or negedge net_w[469]) begin
	#1.26183 net_r[469] <= net_w[469];
end
always @(posedge net_w[470] or negedge net_w[470]) begin
	#5.67823 net_r[470] <= net_w[470];
end
always @(posedge net_w[471] or negedge net_w[471]) begin
	#2.83912 net_r[471] <= net_w[471];
end
always @(posedge net_w[472] or negedge net_w[472]) begin
	#7.57098 net_r[472] <= net_w[472];
end
always @(posedge net_w[473] or negedge net_w[473]) begin
	#2.10305 net_r[473] <= net_w[473];
end
always @(posedge net_w[474] or negedge net_w[474]) begin
	#4.2061 net_r[474] <= net_w[474];
end
always @(posedge net_w[475] or negedge net_w[475]) begin
	#2.94427 net_r[475] <= net_w[475];
end
always @(posedge net_w[476] or negedge net_w[476]) begin
	#2.62881 net_r[476] <= net_w[476];
end
always @(posedge net_w[477] or negedge net_w[477]) begin
	#2.31335 net_r[477] <= net_w[477];
end
always @(posedge net_w[478] or negedge net_w[478]) begin
	#2.83912 net_r[478] <= net_w[478];
end
always @(posedge net_w[479] or negedge net_w[479]) begin
	#1.57729 net_r[479] <= net_w[479];
end
always @(posedge net_w[480] or negedge net_w[480]) begin
	#0.946372 net_r[480] <= net_w[480];
end
always @(posedge net_w[481] or negedge net_w[481]) begin
	#1.9979 net_r[481] <= net_w[481];
end
always @(posedge net_w[482] or negedge net_w[482]) begin
	#1.05152 net_r[482] <= net_w[482];
end
always @(posedge net_w[483] or negedge net_w[483]) begin
	#2.31335 net_r[483] <= net_w[483];
end
always @(posedge net_w[484] or negedge net_w[484]) begin
	#0.525762 net_r[484] <= net_w[484];
end
always @(posedge net_w[485] or negedge net_w[485]) begin
	#1.89274 net_r[485] <= net_w[485];
end
always @(posedge net_w[486] or negedge net_w[486]) begin
	#0.525762 net_r[486] <= net_w[486];
end
always @(posedge net_w[487] or negedge net_w[487]) begin
	#1.47213 net_r[487] <= net_w[487];
end
always @(posedge net_w[488] or negedge net_w[488]) begin
	#0.84122 net_r[488] <= net_w[488];
end
always @(posedge net_w[489] or negedge net_w[489]) begin
	#3.57518 net_r[489] <= net_w[489];
end
always @(posedge net_w[490] or negedge net_w[490]) begin
	#3.99579 net_r[490] <= net_w[490];
end
always @(posedge net_w[491] or negedge net_w[491]) begin
	#3.99579 net_r[491] <= net_w[491];
end
always @(posedge net_w[492] or negedge net_w[492]) begin
	#3.04942 net_r[492] <= net_w[492];
end
always @(posedge net_w[493] or negedge net_w[493]) begin
	#5.04732 net_r[493] <= net_w[493];
end
always @(posedge net_w[494] or negedge net_w[494]) begin
	#5.15247 net_r[494] <= net_w[494];
end
always @(posedge net_w[495] or negedge net_w[495]) begin
	#5.88854 net_r[495] <= net_w[495];
end
always @(posedge net_w[496] or negedge net_w[496]) begin
	#5.36278 net_r[496] <= net_w[496];
end
always @(posedge net_w[497] or negedge net_w[497]) begin
	#3.78549 net_r[497] <= net_w[497];
end
always @(posedge net_w[498] or negedge net_w[498]) begin
	#3.15457 net_r[498] <= net_w[498];
end
always @(posedge net_w[499] or negedge net_w[499]) begin
	#1.68244 net_r[499] <= net_w[499];
end
always @(posedge net_w[500] or negedge net_w[500]) begin
	#1.26183 net_r[500] <= net_w[500];
end
always @(posedge net_w[501] or negedge net_w[501]) begin
	#2.73396 net_r[501] <= net_w[501];
end
always @(posedge net_w[502] or negedge net_w[502]) begin
	#1.26183 net_r[502] <= net_w[502];
end
always @(posedge net_w[503] or negedge net_w[503]) begin
	#1.89274 net_r[503] <= net_w[503];
end
always @(posedge net_w[504] or negedge net_w[504]) begin
	#0.630915 net_r[504] <= net_w[504];
end
always @(posedge net_w[505] or negedge net_w[505]) begin
	#2.31335 net_r[505] <= net_w[505];
end
always @(posedge net_w[506] or negedge net_w[506]) begin
	#1.9979 net_r[506] <= net_w[506];
end
always @(posedge net_w[507] or negedge net_w[507]) begin
	#3.99579 net_r[507] <= net_w[507];
end
always @(posedge net_w[508] or negedge net_w[508]) begin
	#4.2061 net_r[508] <= net_w[508];
end
always @(posedge net_w[509] or negedge net_w[509]) begin
	#5.57308 net_r[509] <= net_w[509];
end
always @(posedge net_w[510] or negedge net_w[510]) begin
	#5.04732 net_r[510] <= net_w[510];
end
always @(posedge net_w[511] or negedge net_w[511]) begin
	#5.78339 net_r[511] <= net_w[511];
end
always @(posedge net_w[512] or negedge net_w[512]) begin
	#4.4164 net_r[512] <= net_w[512];
end
always @(posedge net_w[513] or negedge net_w[513]) begin
	#5.15247 net_r[513] <= net_w[513];
end
always @(posedge net_w[514] or negedge net_w[514]) begin
	#4.52156 net_r[514] <= net_w[514];
end
always @(posedge net_w[515] or negedge net_w[515]) begin
	#1.57729 net_r[515] <= net_w[515];
end
always @(posedge net_w[516] or negedge net_w[516]) begin
	#2.52366 net_r[516] <= net_w[516];
end
always @(posedge net_w[517] or negedge net_w[517]) begin
	#1.47213 net_r[517] <= net_w[517];
end
always @(posedge net_w[518] or negedge net_w[518]) begin
	#2.52366 net_r[518] <= net_w[518];
end
always @(posedge net_w[519] or negedge net_w[519]) begin
	#2.62881 net_r[519] <= net_w[519];
end
always @(posedge net_w[520] or negedge net_w[520]) begin
	#1.57729 net_r[520] <= net_w[520];
end
always @(posedge net_w[521] or negedge net_w[521]) begin
	#2.94427 net_r[521] <= net_w[521];
end
always @(posedge net_w[522] or negedge net_w[522]) begin
	#1.47213 net_r[522] <= net_w[522];
end
always @(posedge net_w[523] or negedge net_w[523]) begin
	#3.36488 net_r[523] <= net_w[523];
end
always @(posedge net_w[524] or negedge net_w[524]) begin
	#1.47213 net_r[524] <= net_w[524];
end
always @(posedge net_w[525] or negedge net_w[525]) begin
	#3.47003 net_r[525] <= net_w[525];
end
always @(posedge net_w[526] or negedge net_w[526]) begin
	#1.47213 net_r[526] <= net_w[526];
end
always @(posedge net_w[527] or negedge net_w[527]) begin
	#1.47213 net_r[527] <= net_w[527];
end
always @(posedge net_w[528] or negedge net_w[528]) begin
	#1.36698 net_r[528] <= net_w[528];
end
always @(posedge net_w[529] or negedge net_w[529]) begin
	#2.10305 net_r[529] <= net_w[529];
end
always @(posedge net_w[530] or negedge net_w[530]) begin
	#1.89274 net_r[530] <= net_w[530];
end
always @(posedge net_w[531] or negedge net_w[531]) begin
	#2.83912 net_r[531] <= net_w[531];
end
always @(posedge net_w[532] or negedge net_w[532]) begin
	#1.89274 net_r[532] <= net_w[532];
end
always @(posedge net_w[533] or negedge net_w[533]) begin
	#2.83912 net_r[533] <= net_w[533];
end
always @(posedge net_w[534] or negedge net_w[534]) begin
	#1.68244 net_r[534] <= net_w[534];
end
always @(posedge net_w[535] or negedge net_w[535]) begin
	#1.89274 net_r[535] <= net_w[535];
end
always @(posedge net_w[536] or negedge net_w[536]) begin
	#2.73396 net_r[536] <= net_w[536];
end
always @(posedge net_w[537] or negedge net_w[537]) begin
	#0.84122 net_r[537] <= net_w[537];
end
always @(posedge net_w[538] or negedge net_w[538]) begin
	#4.83701 net_r[538] <= net_w[538];
end
always @(posedge net_w[539] or negedge net_w[539]) begin
	#1.9979 net_r[539] <= net_w[539];
end
always @(posedge net_w[540] or negedge net_w[540]) begin
	#3.04942 net_r[540] <= net_w[540];
end
always @(posedge net_w[541] or negedge net_w[541]) begin
	#0.630915 net_r[541] <= net_w[541];
end
always @(posedge net_w[542] or negedge net_w[542]) begin
	#2.52366 net_r[542] <= net_w[542];
end
always @(posedge net_w[543] or negedge net_w[543]) begin
	#1.47213 net_r[543] <= net_w[543];
end
always @(posedge net_w[544] or negedge net_w[544]) begin
	#0.525762 net_r[544] <= net_w[544];
end
always @(posedge net_w[545] or negedge net_w[545]) begin
	#1.9979 net_r[545] <= net_w[545];
end
always @(posedge net_w[546] or negedge net_w[546]) begin
	#0.736067 net_r[546] <= net_w[546];
end
always @(posedge net_w[547] or negedge net_w[547]) begin
	#3.68034 net_r[547] <= net_w[547];
end
always @(posedge net_w[548] or negedge net_w[548]) begin
	#3.36488 net_r[548] <= net_w[548];
end
always @(posedge net_w[549] or negedge net_w[549]) begin
	#4.62671 net_r[549] <= net_w[549];
end
always @(posedge net_w[550] or negedge net_w[550]) begin
	#3.47003 net_r[550] <= net_w[550];
end
always @(posedge net_w[551] or negedge net_w[551]) begin
	#2.41851 net_r[551] <= net_w[551];
end
always @(posedge net_w[552] or negedge net_w[552]) begin
	#1.57729 net_r[552] <= net_w[552];
end
always @(posedge net_w[553] or negedge net_w[553]) begin
	#0.84122 net_r[553] <= net_w[553];
end
always @(posedge net_w[554] or negedge net_w[554]) begin
	#4.94217 net_r[554] <= net_w[554];
end
always @(posedge net_w[555] or negedge net_w[555]) begin
	#2.31335 net_r[555] <= net_w[555];
end
always @(posedge net_w[556] or negedge net_w[556]) begin
	#6.62461 net_r[556] <= net_w[556];
end
always @(posedge net_w[557] or negedge net_w[557]) begin
	#2.73396 net_r[557] <= net_w[557];
end
always @(posedge net_w[558] or negedge net_w[558]) begin
	#8.51735 net_r[558] <= net_w[558];
end
always @(posedge net_w[559] or negedge net_w[559]) begin
	#5.99369 net_r[559] <= net_w[559];
end
always @(posedge net_w[560] or negedge net_w[560]) begin
	#2.31335 net_r[560] <= net_w[560];
end
always @(posedge net_w[561] or negedge net_w[561]) begin
	#2.62881 net_r[561] <= net_w[561];
end
always @(posedge net_w[562] or negedge net_w[562]) begin
	#3.04942 net_r[562] <= net_w[562];
end
always @(posedge net_w[563] or negedge net_w[563]) begin
	#1.15668 net_r[563] <= net_w[563];
end
always @(posedge net_w[564] or negedge net_w[564]) begin
	#0.736067 net_r[564] <= net_w[564];
end
always @(posedge net_w[565] or negedge net_w[565]) begin
	#0.946372 net_r[565] <= net_w[565];
end
always @(posedge net_w[566] or negedge net_w[566]) begin
	#0.736067 net_r[566] <= net_w[566];
end
always @(posedge net_w[567] or negedge net_w[567]) begin
	#0.946372 net_r[567] <= net_w[567];
end
always @(posedge net_w[568] or negedge net_w[568]) begin
	#0.736067 net_r[568] <= net_w[568];
end
always @(posedge net_w[569] or negedge net_w[569]) begin
	#0.946372 net_r[569] <= net_w[569];
end
always @(posedge net_w[570] or negedge net_w[570]) begin
	#0.736067 net_r[570] <= net_w[570];
end
always @(posedge net_w[571] or negedge net_w[571]) begin
	#0.946372 net_r[571] <= net_w[571];
end
always @(posedge net_w[572] or negedge net_w[572]) begin
	#0.736067 net_r[572] <= net_w[572];
end
always @(posedge net_w[573] or negedge net_w[573]) begin
	#0.946372 net_r[573] <= net_w[573];
end
always @(posedge net_w[574] or negedge net_w[574]) begin
	#0.736067 net_r[574] <= net_w[574];
end
always @(posedge net_w[575] or negedge net_w[575]) begin
	#0.946372 net_r[575] <= net_w[575];
end
always @(posedge net_w[576] or negedge net_w[576]) begin
	#0.736067 net_r[576] <= net_w[576];
end
always @(posedge net_w[577] or negedge net_w[577]) begin
	#0.946372 net_r[577] <= net_w[577];
end
always @(posedge net_w[578] or negedge net_w[578]) begin
	#0.736067 net_r[578] <= net_w[578];
end
always @(posedge net_w[579] or negedge net_w[579]) begin
	#1.47213 net_r[579] <= net_w[579];
end
always @(posedge net_w[580] or negedge net_w[580]) begin
	#1.47213 net_r[580] <= net_w[580];
end
always @(posedge net_w[581] or negedge net_w[581]) begin
	#1.47213 net_r[581] <= net_w[581];
end
always @(posedge net_w[582] or negedge net_w[582]) begin
	#1.47213 net_r[582] <= net_w[582];
end
always @(posedge net_w[583] or negedge net_w[583]) begin
	#1.68244 net_r[583] <= net_w[583];
end
always @(posedge net_w[584] or negedge net_w[584]) begin
	#1.26183 net_r[584] <= net_w[584];
end
always @(posedge net_w[585] or negedge net_w[585]) begin
	#1.47213 net_r[585] <= net_w[585];
end
always @(posedge net_w[586] or negedge net_w[586]) begin
	#1.47213 net_r[586] <= net_w[586];
end
always @(posedge net_w[587] or negedge net_w[587]) begin
	#3.15457 net_r[587] <= net_w[587];
end
always @(posedge net_w[588] or negedge net_w[588]) begin
	#2.52366 net_r[588] <= net_w[588];
end
always @(posedge net_w[589] or negedge net_w[589]) begin
	#2.73396 net_r[589] <= net_w[589];
end
always @(posedge net_w[590] or negedge net_w[590]) begin
	#2.52366 net_r[590] <= net_w[590];
end
always @(posedge net_w[591] or negedge net_w[591]) begin
	#5.88854 net_r[591] <= net_w[591];
end
always @(posedge net_w[592] or negedge net_w[592]) begin
	#4.62671 net_r[592] <= net_w[592];
end
always @(posedge net_w[593] or negedge net_w[593]) begin
	#0.946372 net_r[593] <= net_w[593];
end
always @(posedge net_w[594] or negedge net_w[594]) begin
	#0.736067 net_r[594] <= net_w[594];
end
always @(posedge net_w[595] or negedge net_w[595]) begin
	#0.946372 net_r[595] <= net_w[595];
end
always @(posedge net_w[596] or negedge net_w[596]) begin
	#0.84122 net_r[596] <= net_w[596];
end
always @(posedge net_w[597] or negedge net_w[597]) begin
	#0.946372 net_r[597] <= net_w[597];
end
always @(posedge net_w[598] or negedge net_w[598]) begin
	#0.736067 net_r[598] <= net_w[598];
end
always @(posedge net_w[599] or negedge net_w[599]) begin
	#0.946372 net_r[599] <= net_w[599];
end
always @(posedge net_w[600] or negedge net_w[600]) begin
	#1.26183 net_r[600] <= net_w[600];
end
always @(posedge net_w[601] or negedge net_w[601]) begin
	#0.946372 net_r[601] <= net_w[601];
end
always @(posedge net_w[602] or negedge net_w[602]) begin
	#1.26183 net_r[602] <= net_w[602];
end
always @(posedge net_w[603] or negedge net_w[603]) begin
	#0.946372 net_r[603] <= net_w[603];
end
always @(posedge net_w[604] or negedge net_w[604]) begin
	#1.89274 net_r[604] <= net_w[604];
end
always @(posedge net_w[605] or negedge net_w[605]) begin
	#0.946372 net_r[605] <= net_w[605];
end
always @(posedge net_w[606] or negedge net_w[606]) begin
	#1.26183 net_r[606] <= net_w[606];
end
always @(posedge net_w[607] or negedge net_w[607]) begin
	#7.67613 net_r[607] <= net_w[607];
end
always @(posedge net_w[608] or negedge net_w[608]) begin
	#2.94427 net_r[608] <= net_w[608];
end
always @(posedge net_w[609] or negedge net_w[609]) begin
	#1.47213 net_r[609] <= net_w[609];
end
always @(posedge net_w[610] or negedge net_w[610]) begin
	#1.68244 net_r[610] <= net_w[610];
end
always @(posedge net_w[611] or negedge net_w[611]) begin
	#1.57729 net_r[611] <= net_w[611];
end
always @(posedge net_w[612] or negedge net_w[612]) begin
	#1.36698 net_r[612] <= net_w[612];
end
always @(posedge net_w[613] or negedge net_w[613]) begin
	#0.84122 net_r[613] <= net_w[613];
end
always @(posedge net_w[614] or negedge net_w[614]) begin
	#1.57729 net_r[614] <= net_w[614];
end
always @(posedge net_w[615] or negedge net_w[615]) begin
	#1.26183 net_r[615] <= net_w[615];
end
always @(posedge net_w[616] or negedge net_w[616]) begin
	#2.83912 net_r[616] <= net_w[616];
end
always @(posedge net_w[617] or negedge net_w[617]) begin
	#2.52366 net_r[617] <= net_w[617];
end
always @(posedge net_w[618] or negedge net_w[618]) begin
	#2.62881 net_r[618] <= net_w[618];
end
always @(posedge net_w[619] or negedge net_w[619]) begin
	#2.31335 net_r[619] <= net_w[619];
end
always @(posedge net_w[620] or negedge net_w[620]) begin
	#5.04732 net_r[620] <= net_w[620];
end
always @(posedge net_w[621] or negedge net_w[621]) begin
	#3.99579 net_r[621] <= net_w[621];
end
always @(posedge net_w[622] or negedge net_w[622]) begin
	#1.68244 net_r[622] <= net_w[622];
end
always @(posedge net_w[623] or negedge net_w[623]) begin
	#0.84122 net_r[623] <= net_w[623];
end
always @(posedge net_w[624] or negedge net_w[624]) begin
	#1.05152 net_r[624] <= net_w[624];
end
always @(posedge net_w[625] or negedge net_w[625]) begin
	#0.736067 net_r[625] <= net_w[625];
end
always @(posedge net_w[626] or negedge net_w[626]) begin
	#1.26183 net_r[626] <= net_w[626];
end
always @(posedge net_w[627] or negedge net_w[627]) begin
	#0.736067 net_r[627] <= net_w[627];
end
always @(posedge net_w[628] or negedge net_w[628]) begin
	#1.05152 net_r[628] <= net_w[628];
end
always @(posedge net_w[629] or negedge net_w[629]) begin
	#2.62881 net_r[629] <= net_w[629];
end
always @(posedge net_w[630] or negedge net_w[630]) begin
	#1.05152 net_r[630] <= net_w[630];
end
always @(posedge net_w[631] or negedge net_w[631]) begin
	#1.47213 net_r[631] <= net_w[631];
end
always @(posedge net_w[632] or negedge net_w[632]) begin
	#0.946372 net_r[632] <= net_w[632];
end
always @(posedge net_w[633] or negedge net_w[633]) begin
	#1.36698 net_r[633] <= net_w[633];
end
always @(posedge net_w[634] or negedge net_w[634]) begin
	#7.78128 net_r[634] <= net_w[634];
end
always @(posedge net_w[635] or negedge net_w[635]) begin
	#1.78759 net_r[635] <= net_w[635];
end
always @(posedge net_w[636] or negedge net_w[636]) begin
	#1.68244 net_r[636] <= net_w[636];
end
always @(posedge net_w[637] or negedge net_w[637]) begin
	#1.78759 net_r[637] <= net_w[637];
end
always @(posedge net_w[638] or negedge net_w[638]) begin
	#2.83912 net_r[638] <= net_w[638];
end
always @(posedge net_w[639] or negedge net_w[639]) begin
	#1.47213 net_r[639] <= net_w[639];
end
always @(posedge net_w[640] or negedge net_w[640]) begin
	#1.36698 net_r[640] <= net_w[640];
end
always @(posedge net_w[641] or negedge net_w[641]) begin
	#6.94006 net_r[641] <= net_w[641];
end
always @(posedge net_w[642] or negedge net_w[642]) begin
	#3.25973 net_r[642] <= net_w[642];
end
always @(posedge net_w[643] or negedge net_w[643]) begin
	#3.25973 net_r[643] <= net_w[643];
end
always @(posedge net_w[644] or negedge net_w[644]) begin
	#2.31335 net_r[644] <= net_w[644];
end
always @(posedge net_w[645] or negedge net_w[645]) begin
	#1.57729 net_r[645] <= net_w[645];
end
always @(posedge net_w[646] or negedge net_w[646]) begin
	#4.52156 net_r[646] <= net_w[646];
end
always @(posedge net_w[647] or negedge net_w[647]) begin
	#2.62881 net_r[647] <= net_w[647];
end
always @(posedge net_w[648] or negedge net_w[648]) begin
	#1.05152 net_r[648] <= net_w[648];
end
always @(posedge net_w[649] or negedge net_w[649]) begin
	#0.84122 net_r[649] <= net_w[649];
end
always @(posedge net_w[650] or negedge net_w[650]) begin
	#1.15668 net_r[650] <= net_w[650];
end
always @(posedge net_w[651] or negedge net_w[651]) begin
	#0.84122 net_r[651] <= net_w[651];
end
always @(posedge net_w[652] or negedge net_w[652]) begin
	#1.68244 net_r[652] <= net_w[652];
end
always @(posedge net_w[653] or negedge net_w[653]) begin
	#1.57729 net_r[653] <= net_w[653];
end
always @(posedge net_w[654] or negedge net_w[654]) begin
	#1.05152 net_r[654] <= net_w[654];
end
always @(posedge net_w[655] or negedge net_w[655]) begin
	#0.84122 net_r[655] <= net_w[655];
end
always @(posedge net_w[656] or negedge net_w[656]) begin
	#1.36698 net_r[656] <= net_w[656];
end
always @(posedge net_w[657] or negedge net_w[657]) begin
	#0.84122 net_r[657] <= net_w[657];
end
always @(posedge net_w[658] or negedge net_w[658]) begin
	#1.05152 net_r[658] <= net_w[658];
end
always @(posedge net_w[659] or negedge net_w[659]) begin
	#0.84122 net_r[659] <= net_w[659];
end
always @(posedge net_w[660] or negedge net_w[660]) begin
	#1.68244 net_r[660] <= net_w[660];
end
always @(posedge net_w[661] or negedge net_w[661]) begin
	#2.2082 net_r[661] <= net_w[661];
end
always @(posedge net_w[662] or negedge net_w[662]) begin
	#2.62881 net_r[662] <= net_w[662];
end
always @(posedge net_w[663] or negedge net_w[663]) begin
	#1.47213 net_r[663] <= net_w[663];
end
always @(posedge net_w[664] or negedge net_w[664]) begin
	#1.89274 net_r[664] <= net_w[664];
end
always @(posedge net_w[665] or negedge net_w[665]) begin
	#1.68244 net_r[665] <= net_w[665];
end
always @(posedge net_w[666] or negedge net_w[666]) begin
	#4.31125 net_r[666] <= net_w[666];
end
always @(posedge net_w[667] or negedge net_w[667]) begin
	#4.10095 net_r[667] <= net_w[667];
end
always @(posedge net_w[668] or negedge net_w[668]) begin
	#6.72976 net_r[668] <= net_w[668];
end
always @(posedge net_w[669] or negedge net_w[669]) begin
	#2.10305 net_r[669] <= net_w[669];
end
always @(posedge net_w[670] or negedge net_w[670]) begin
	#1.68244 net_r[670] <= net_w[670];
end
always @(posedge net_w[671] or negedge net_w[671]) begin
	#1.15668 net_r[671] <= net_w[671];
end
always @(posedge net_w[672] or negedge net_w[672]) begin
	#0.84122 net_r[672] <= net_w[672];
end
always @(posedge net_w[673] or negedge net_w[673]) begin
	#1.26183 net_r[673] <= net_w[673];
end
always @(posedge net_w[674] or negedge net_w[674]) begin
	#0.946372 net_r[674] <= net_w[674];
end
always @(posedge net_w[675] or negedge net_w[675]) begin
	#2.41851 net_r[675] <= net_w[675];
end
always @(posedge net_w[676] or negedge net_w[676]) begin
	#0.84122 net_r[676] <= net_w[676];
end
always @(posedge net_w[677] or negedge net_w[677]) begin
	#1.57729 net_r[677] <= net_w[677];
end
always @(posedge net_w[678] or negedge net_w[678]) begin
	#2.52366 net_r[678] <= net_w[678];
end
always @(posedge net_w[679] or negedge net_w[679]) begin
	#1.05152 net_r[679] <= net_w[679];
end
always @(posedge net_w[680] or negedge net_w[680]) begin
	#1.78759 net_r[680] <= net_w[680];
end
always @(posedge net_w[681] or negedge net_w[681]) begin
	#6.204 net_r[681] <= net_w[681];
end
always @(posedge net_w[682] or negedge net_w[682]) begin
	#2.2082 net_r[682] <= net_w[682];
end
always @(posedge net_w[683] or negedge net_w[683]) begin
	#4.2061 net_r[683] <= net_w[683];
end
always @(posedge net_w[684] or negedge net_w[684]) begin
	#1.9979 net_r[684] <= net_w[684];
end
always @(posedge net_w[685] or negedge net_w[685]) begin
	#0.84122 net_r[685] <= net_w[685];
end
always @(posedge net_w[686] or negedge net_w[686]) begin
	#1.78759 net_r[686] <= net_w[686];
end
always @(posedge net_w[687] or negedge net_w[687]) begin
	#1.57729 net_r[687] <= net_w[687];
end
always @(posedge net_w[688] or negedge net_w[688]) begin
	#4.52156 net_r[688] <= net_w[688];
end
always @(posedge net_w[689] or negedge net_w[689]) begin
	#4.52156 net_r[689] <= net_w[689];
end
always @(posedge net_w[690] or negedge net_w[690]) begin
	#5.36278 net_r[690] <= net_w[690];
end
always @(posedge net_w[691] or negedge net_w[691]) begin
	#1.78759 net_r[691] <= net_w[691];
end
always @(posedge net_w[692] or negedge net_w[692]) begin
	#0.84122 net_r[692] <= net_w[692];
end
always @(posedge net_w[693] or negedge net_w[693]) begin
	#1.15668 net_r[693] <= net_w[693];
end
always @(posedge net_w[694] or negedge net_w[694]) begin
	#0.946372 net_r[694] <= net_w[694];
end
always @(posedge net_w[695] or negedge net_w[695]) begin
	#1.15668 net_r[695] <= net_w[695];
end
always @(posedge net_w[696] or negedge net_w[696]) begin
	#7.57098 net_r[696] <= net_w[696];
end
always @(posedge net_w[697] or negedge net_w[697]) begin
	#1.89274 net_r[697] <= net_w[697];
end
always @(posedge net_w[698] or negedge net_w[698]) begin
	#1.68244 net_r[698] <= net_w[698];
end
always @(posedge net_w[699] or negedge net_w[699]) begin
	#1.15668 net_r[699] <= net_w[699];
end
always @(posedge net_w[700] or negedge net_w[700]) begin
	#0.946372 net_r[700] <= net_w[700];
end
always @(posedge net_w[701] or negedge net_w[701]) begin
	#1.15668 net_r[701] <= net_w[701];
end
always @(posedge net_w[702] or negedge net_w[702]) begin
	#0.946372 net_r[702] <= net_w[702];
end
always @(posedge net_w[703] or negedge net_w[703]) begin
	#1.89274 net_r[703] <= net_w[703];
end
always @(posedge net_w[704] or negedge net_w[704]) begin
	#2.10305 net_r[704] <= net_w[704];
end
always @(posedge net_w[705] or negedge net_w[705]) begin
	#1.15668 net_r[705] <= net_w[705];
end
always @(posedge net_w[706] or negedge net_w[706]) begin
	#2.62881 net_r[706] <= net_w[706];
end
always @(posedge net_w[707] or negedge net_w[707]) begin
	#7.36067 net_r[707] <= net_w[707];
end
always @(posedge net_w[708] or negedge net_w[708]) begin
	#2.83912 net_r[708] <= net_w[708];
end
always @(posedge net_w[709] or negedge net_w[709]) begin
	#9.14826 net_r[709] <= net_w[709];
end
always @(posedge net_w[710] or negedge net_w[710]) begin
	#4.10095 net_r[710] <= net_w[710];
end
always @(posedge net_w[711] or negedge net_w[711]) begin
	#7.04522 net_r[711] <= net_w[711];
end
always @(posedge net_w[712] or negedge net_w[712]) begin
	#0.946372 net_r[712] <= net_w[712];
end
always @(posedge net_w[713] or negedge net_w[713]) begin
	#1.26183 net_r[713] <= net_w[713];
end
always @(posedge net_w[714] or negedge net_w[714]) begin
	#0.946372 net_r[714] <= net_w[714];
end
always @(posedge net_w[715] or negedge net_w[715]) begin
	#4.62671 net_r[715] <= net_w[715];
end
always @(posedge net_w[716] or negedge net_w[716]) begin
	#1.05152 net_r[716] <= net_w[716];
end
always @(posedge net_w[717] or negedge net_w[717]) begin
	#2.41851 net_r[717] <= net_w[717];
end
always @(posedge net_w[718] or negedge net_w[718]) begin
	#1.78759 net_r[718] <= net_w[718];
end
always @(posedge net_w[719] or negedge net_w[719]) begin
	#1.26183 net_r[719] <= net_w[719];
end
always @(posedge net_w[720] or negedge net_w[720]) begin
	#2.83912 net_r[720] <= net_w[720];
end
always @(posedge net_w[721] or negedge net_w[721]) begin
	#4.62671 net_r[721] <= net_w[721];
end
always @(posedge net_w[722] or negedge net_w[722]) begin
	#2.2082 net_r[722] <= net_w[722];
end
always @(posedge net_w[723] or negedge net_w[723]) begin
	#5.46793 net_r[723] <= net_w[723];
end
always @(posedge net_w[724] or negedge net_w[724]) begin
	#1.15668 net_r[724] <= net_w[724];
end
always @(posedge net_w[725] or negedge net_w[725]) begin
	#1.78759 net_r[725] <= net_w[725];
end
always @(posedge net_w[726] or negedge net_w[726]) begin
	#5.46793 net_r[726] <= net_w[726];
end
always @(posedge net_w[727] or negedge net_w[727]) begin
	#4.2061 net_r[727] <= net_w[727];
end
always @(posedge net_w[728] or negedge net_w[728]) begin
	#2.62881 net_r[728] <= net_w[728];
end
always @(posedge net_w[729] or negedge net_w[729]) begin
	#7.57098 net_r[729] <= net_w[729];
end
always @(posedge net_w[730] or negedge net_w[730]) begin
	#1.26183 net_r[730] <= net_w[730];
end
always @(posedge net_w[731] or negedge net_w[731]) begin
	#0.946372 net_r[731] <= net_w[731];
end
always @(posedge net_w[732] or negedge net_w[732]) begin
	#1.47213 net_r[732] <= net_w[732];
end
always @(posedge net_w[733] or negedge net_w[733]) begin
	#1.26183 net_r[733] <= net_w[733];
end
always @(posedge net_w[734] or negedge net_w[734]) begin
	#3.15457 net_r[734] <= net_w[734];
end
always @(posedge net_w[735] or negedge net_w[735]) begin
	#2.31335 net_r[735] <= net_w[735];
end
always @(posedge net_w[736] or negedge net_w[736]) begin
	#1.47213 net_r[736] <= net_w[736];
end
always @(posedge net_w[737] or negedge net_w[737]) begin
	#2.31335 net_r[737] <= net_w[737];
end
always @(posedge net_w[738] or negedge net_w[738]) begin
	#6.30915 net_r[738] <= net_w[738];
end
always @(posedge net_w[739] or negedge net_w[739]) begin
	#2.73396 net_r[739] <= net_w[739];
end
always @(posedge net_w[740] or negedge net_w[740]) begin
	#5.67823 net_r[740] <= net_w[740];
end
always @(posedge net_w[741] or negedge net_w[741]) begin
	#1.47213 net_r[741] <= net_w[741];
end
always @(posedge net_w[742] or negedge net_w[742]) begin
	#1.26183 net_r[742] <= net_w[742];
end
always @(posedge net_w[743] or negedge net_w[743]) begin
	#6.94006 net_r[743] <= net_w[743];
end
always @(posedge net_w[744] or negedge net_w[744]) begin
	#3.36488 net_r[744] <= net_w[744];
end
always @(posedge net_w[745] or negedge net_w[745]) begin
	#5.67823 net_r[745] <= net_w[745];
end
always @(posedge net_w[746] or negedge net_w[746]) begin
	#1.36698 net_r[746] <= net_w[746];
end
always @(posedge net_w[747] or negedge net_w[747]) begin
	#1.26183 net_r[747] <= net_w[747];
end
always @(posedge net_w[748] or negedge net_w[748]) begin
	#1.36698 net_r[748] <= net_w[748];
end
always @(posedge net_w[749] or negedge net_w[749]) begin
	#1.26183 net_r[749] <= net_w[749];
end
always @(posedge net_w[750] or negedge net_w[750]) begin
	#1.36698 net_r[750] <= net_w[750];
end
always @(posedge net_w[751] or negedge net_w[751]) begin
	#1.15668 net_r[751] <= net_w[751];
end
always @(posedge net_w[752] or negedge net_w[752]) begin
	#1.47213 net_r[752] <= net_w[752];
end
always @(posedge net_w[753] or negedge net_w[753]) begin
	#1.15668 net_r[753] <= net_w[753];
end
always @(posedge net_w[754] or negedge net_w[754]) begin
	#2.83912 net_r[754] <= net_w[754];
end
always @(posedge net_w[755] or negedge net_w[755]) begin
	#3.15457 net_r[755] <= net_w[755];
end
always @(posedge net_w[756] or negedge net_w[756]) begin
	#2.62881 net_r[756] <= net_w[756];
end
always @(posedge net_w[757] or negedge net_w[757]) begin
	#2.41851 net_r[757] <= net_w[757];
end
always @(posedge net_w[758] or negedge net_w[758]) begin
	#6.204 net_r[758] <= net_w[758];
end
always @(posedge net_w[759] or negedge net_w[759]) begin
	#5.25762 net_r[759] <= net_w[759];
end
always @(posedge net_w[760] or negedge net_w[760]) begin
	#4.31125 net_r[760] <= net_w[760];
end
always @(posedge net_w[761] or negedge net_w[761]) begin
	#1.47213 net_r[761] <= net_w[761];
end
always @(posedge net_w[762] or negedge net_w[762]) begin
	#1.26183 net_r[762] <= net_w[762];
end
always @(posedge net_w[763] or negedge net_w[763]) begin
	#1.47213 net_r[763] <= net_w[763];
end
always @(posedge net_w[764] or negedge net_w[764]) begin
	#2.31335 net_r[764] <= net_w[764];
end
always @(posedge net_w[765] or negedge net_w[765]) begin
	#1.47213 net_r[765] <= net_w[765];
end
always @(posedge net_w[766] or negedge net_w[766]) begin
	#2.31335 net_r[766] <= net_w[766];
end
always @(posedge net_w[767] or negedge net_w[767]) begin
	#5.88854 net_r[767] <= net_w[767];
end
always @(posedge net_w[768] or negedge net_w[768]) begin
	#2.52366 net_r[768] <= net_w[768];
end
always @(posedge net_w[769] or negedge net_w[769]) begin
	#3.57518 net_r[769] <= net_w[769];
end
always @(posedge net_w[770] or negedge net_w[770]) begin
	#1.47213 net_r[770] <= net_w[770];
end
always @(posedge net_w[771] or negedge net_w[771]) begin
	#1.26183 net_r[771] <= net_w[771];
end
always @(posedge net_w[772] or negedge net_w[772]) begin
	#4.83701 net_r[772] <= net_w[772];
end
always @(posedge net_w[773] or negedge net_w[773]) begin
	#3.57518 net_r[773] <= net_w[773];
end
always @(posedge net_w[774] or negedge net_w[774]) begin
	#3.57518 net_r[774] <= net_w[774];
end
always @(posedge net_w[775] or negedge net_w[775]) begin
	#1.68244 net_r[775] <= net_w[775];
end
always @(posedge net_w[776] or negedge net_w[776]) begin
	#1.36698 net_r[776] <= net_w[776];
end
always @(posedge net_w[777] or negedge net_w[777]) begin
	#1.68244 net_r[777] <= net_w[777];
end
always @(posedge net_w[778] or negedge net_w[778]) begin
	#2.62881 net_r[778] <= net_w[778];
end
always @(posedge net_w[779] or negedge net_w[779]) begin
	#2.83912 net_r[779] <= net_w[779];
end
always @(posedge net_w[780] or negedge net_w[780]) begin
	#3.99579 net_r[780] <= net_w[780];
end
always @(posedge net_w[781] or negedge net_w[781]) begin
	#5.25762 net_r[781] <= net_w[781];
end
always @(posedge net_w[782] or negedge net_w[782]) begin
	#4.4164 net_r[782] <= net_w[782];
end
always @(posedge net_w[783] or negedge net_w[783]) begin
	#1.78759 net_r[783] <= net_w[783];
end
always @(posedge net_w[784] or negedge net_w[784]) begin
	#1.47213 net_r[784] <= net_w[784];
end
always @(posedge net_w[785] or negedge net_w[785]) begin
	#2.73396 net_r[785] <= net_w[785];
end
always @(posedge net_w[786] or negedge net_w[786]) begin
	#2.10305 net_r[786] <= net_w[786];
end
always @(posedge net_w[787] or negedge net_w[787]) begin
	#5.25762 net_r[787] <= net_w[787];
end
always @(posedge net_w[788] or negedge net_w[788]) begin
	#2.10305 net_r[788] <= net_w[788];
end
always @(posedge net_w[789] or negedge net_w[789]) begin
	#7.15037 net_r[789] <= net_w[789];
end
always @(posedge net_w[790] or negedge net_w[790]) begin
	#1.89274 net_r[790] <= net_w[790];
end
always @(posedge net_w[791] or negedge net_w[791]) begin
	#4.4164 net_r[791] <= net_w[791];
end
always @(posedge net_w[792] or negedge net_w[792]) begin
	#2.10305 net_r[792] <= net_w[792];
end
always @(posedge net_w[793] or negedge net_w[793]) begin
	#5.88854 net_r[793] <= net_w[793];
end
always @(posedge net_w[794] or negedge net_w[794]) begin
	#5.78339 net_r[794] <= net_w[794];
end
always @(posedge net_w[795] or negedge net_w[795]) begin
	#2.31335 net_r[795] <= net_w[795];
end
always @(posedge net_w[796] or negedge net_w[796]) begin
	#8.09674 net_r[796] <= net_w[796];
end
always @(posedge net_w[797] or negedge net_w[797]) begin
	#2.10305 net_r[797] <= net_w[797];
end
always @(posedge net_w[798] or negedge net_w[798]) begin
	#4.10095 net_r[798] <= net_w[798];
end
always @(posedge net_w[799] or negedge net_w[799]) begin
	#2.31335 net_r[799] <= net_w[799];
end
always @(posedge net_w[800] or negedge net_w[800]) begin
	#9.35857 net_r[800] <= net_w[800];
end
always @(posedge net_w[801] or negedge net_w[801]) begin
	#10.1998 net_r[801] <= net_w[801];
end
always @(posedge net_w[802] or negedge net_w[802]) begin
	#5.36278 net_r[802] <= net_w[802];
end
always @(posedge net_w[803] or negedge net_w[803]) begin
	#4.10095 net_r[803] <= net_w[803];
end
always @(posedge net_w[804] or negedge net_w[804]) begin
	#6.62461 net_r[804] <= net_w[804];
end
always @(posedge net_w[805] or negedge net_w[805]) begin
	#4.10095 net_r[805] <= net_w[805];
end
always @(posedge net_w[806] or negedge net_w[806]) begin
	#3.36488 net_r[806] <= net_w[806];
end
always @(posedge net_w[807] or negedge net_w[807]) begin
	#1.78759 net_r[807] <= net_w[807];
end
always @(posedge net_w[808] or negedge net_w[808]) begin
	#3.36488 net_r[808] <= net_w[808];
end
always @(posedge net_w[809] or negedge net_w[809]) begin
	#2.31335 net_r[809] <= net_w[809];
end
always @(posedge net_w[810] or negedge net_w[810]) begin
	#2.62881 net_r[810] <= net_w[810];
end
always @(posedge net_w[811] or negedge net_w[811]) begin
	#2.41851 net_r[811] <= net_w[811];
end
always @(posedge net_w[812] or negedge net_w[812]) begin
	#3.47003 net_r[812] <= net_w[812];
end
always @(posedge net_w[813] or negedge net_w[813]) begin
	#6.4143 net_r[813] <= net_w[813];
end
always @(posedge net_w[814] or negedge net_w[814]) begin
	#9.04311 net_r[814] <= net_w[814];
end
always @(posedge net_w[815] or negedge net_w[815]) begin
	#10.1998 net_r[815] <= net_w[815];
end
always @(posedge net_w[816] or negedge net_w[816]) begin
	#24.2902 net_r[816] <= net_w[816];
end
always @(posedge net_w[817] or negedge net_w[817]) begin
	#10.0946 net_r[817] <= net_w[817];
end
always @(posedge net_w[818] or negedge net_w[818]) begin
	#9.46372 net_r[818] <= net_w[818];
end
always @(posedge net_w[819] or negedge net_w[819]) begin
	#13.6698 net_r[819] <= net_w[819];
end
always @(posedge net_w[820] or negedge net_w[820]) begin
	#7.04522 net_r[820] <= net_w[820];
end
always @(posedge net_w[821] or negedge net_w[821]) begin
	#9.04311 net_r[821] <= net_w[821];
end
always @(posedge net_w[822] or negedge net_w[822]) begin
	#6.72976 net_r[822] <= net_w[822];
end
always @(posedge net_w[823] or negedge net_w[823]) begin
	#9.35857 net_r[823] <= net_w[823];
end
always @(posedge net_w[824] or negedge net_w[824]) begin
	#8.6225 net_r[824] <= net_w[824];
end
always @(posedge net_w[825] or negedge net_w[825]) begin
	#11.8822 net_r[825] <= net_w[825];
end
always @(posedge net_w[826] or negedge net_w[826]) begin
	#13.2492 net_r[826] <= net_w[826];
end
LSmitll_XORT_v2p1_optimized XOR2T_0 (.a(net_r[248]), .b(net_r[279]), .clk(net_r[333]), .q(net_w[18]));
LSmitll_XORT_v2p1_optimized XOR2T_1 (.a(net_r[310]), .b(net_r[312]), .clk(net_r[364]), .q(net_w[198]));
LSmitll_AND2T AND2T_2 (.a(net_r[249]), .b(net_r[280]), .clk(net_r[335]), .q(net_w[176]));
LSmitll_AND2T AND2T_3 (.a(net_r[311]), .b(net_r[313]), .clk(net_r[366]), .q(net_w[20]));
LSmitll_OR2T_v2p1_optimized OR2T_4 (.a(net_r[19]), .b(net_r[20]), .clk(net_r[395]), .q(net_w[21]));
LSmitll_XORT_v2p1_optimized XOR2T_5 (.a(net_r[250]), .b(net_r[281]), .clk(net_r[367]), .q(net_w[22]));
LSmitll_XORT_v2p1_optimized XOR2T_6 (.a(net_r[314]), .b(net_r[316]), .clk(net_r[421]), .q(net_w[211]));
LSmitll_XORT_v2p1_optimized XOR2T_7 (.a(net_r[252]), .b(net_r[283]), .clk(net_r[396]), .q(net_w[23]));
LSmitll_AND2T AND2T_8 (.a(net_r[251]), .b(net_r[282]), .clk(net_r[369]), .q(net_w[177]));
LSmitll_AND2T AND2T_9 (.a(net_r[315]), .b(net_r[317]), .clk(net_r[423]), .q(net_w[25]));
LSmitll_OR2T_v2p1_optimized OR2T_10 (.a(net_r[24]), .b(net_r[25]), .clk(net_r[424]), .q(net_w[26]));
LSmitll_XORT_v2p1_optimized XOR2T_11 (.a(net_r[318]), .b(net_r[320]), .clk(net_r[446]), .q(net_w[222]));
LSmitll_AND2T AND2T_12 (.a(net_r[253]), .b(net_r[284]), .clk(net_r[398]), .q(net_w[178]));
LSmitll_AND2T AND2T_13 (.a(net_r[319]), .b(net_r[321]), .clk(net_r[448]), .q(net_w[28]));
LSmitll_OR2T_v2p1_optimized OR2T_14 (.a(net_r[27]), .b(net_r[28]), .clk(net_r[470]), .q(net_w[29]));
LSmitll_XORT_v2p1_optimized XOR2T_15 (.a(net_r[256]), .b(net_r[287]), .clk(net_r[447]), .q(net_w[30]));
LSmitll_XORT_v2p1_optimized XOR2T_16 (.a(net_r[30]), .b(net_r[322]), .clk(net_r[489]), .q(net_w[231]));
LSmitll_XORT_v2p1_optimized XOR2T_17 (.a(net_r[261]), .b(net_r[292]), .clk(net_r[471]), .q(net_w[31]));
LSmitll_AND2T AND2T_18 (.a(net_r[257]), .b(net_r[288]), .clk(net_r[451]), .q(net_w[179]));
LSmitll_OR2T_v2p1_optimized OR2T_19 (.a(net_r[258]), .b(net_r[289]), .clk(net_r[449]), .q(net_w[33]));
LSmitll_AND2T AND2T_20 (.a(net_r[33]), .b(net_r[323]), .clk(net_r[491]), .q(net_w[34]));
LSmitll_OR2T_v2p1_optimized OR2T_21 (.a(net_r[32]), .b(net_r[34]), .clk(net_r[492]), .q(net_w[35]));
LSmitll_XORT_v2p1_optimized XOR2T_22 (.a(net_r[31]), .b(net_r[324]), .clk(net_r[509]), .q(net_w[238]));
LSmitll_XORT_v2p1_optimized XOR2T_23 (.a(net_r[266]), .b(net_r[297]), .clk(net_r[493]), .q(net_w[36]));
LSmitll_AND2T AND2T_24 (.a(net_r[262]), .b(net_r[293]), .clk(net_r[474]), .q(net_w[180]));
LSmitll_OR2T_v2p1_optimized OR2T_25 (.a(net_r[263]), .b(net_r[294]), .clk(net_r[473]), .q(net_w[38]));
LSmitll_AND2T AND2T_26 (.a(net_r[38]), .b(net_r[325]), .clk(net_r[511]), .q(net_w[39]));
LSmitll_OR2T_v2p1_optimized OR2T_27 (.a(net_r[37]), .b(net_r[39]), .clk(net_r[525]), .q(net_w[40]));
LSmitll_XORT_v2p1_optimized XOR2T_28 (.a(net_r[36]), .b(net_r[326]), .clk(net_r[540]), .q(net_w[243]));
LSmitll_XORT_v2p1_optimized XOR2T_29 (.a(net_r[271]), .b(net_r[302]), .clk(net_r[510]), .q(net_w[41]));
LSmitll_AND2T AND2T_30 (.a(net_r[267]), .b(net_r[298]), .clk(net_r[496]), .q(net_w[181]));
LSmitll_OR2T_v2p1_optimized OR2T_31 (.a(net_r[268]), .b(net_r[299]), .clk(net_r[495]), .q(net_w[43]));
LSmitll_AND2T AND2T_32 (.a(net_r[43]), .b(net_r[327]), .clk(net_r[542]), .q(net_w[44]));
LSmitll_OR2T_v2p1_optimized OR2T_33 (.a(net_r[42]), .b(net_r[44]), .clk(net_r[541]), .q(net_w[45]));
LSmitll_XORT_v2p1_optimized XOR2T_34 (.a(net_r[41]), .b(net_r[328]), .clk(net_r[550]), .q(net_w[246]));
LSmitll_XORT_v2p1_optimized XOR2T_35 (.a(net_r[276]), .b(net_r[307]), .clk(net_r[526]), .q(net_w[46]));
LSmitll_AND2T AND2T_36 (.a(net_r[272]), .b(net_r[303]), .clk(net_r[514]), .q(net_w[182]));
LSmitll_OR2T_v2p1_optimized OR2T_37 (.a(net_r[273]), .b(net_r[304]), .clk(net_r[512]), .q(net_w[48]));
LSmitll_AND2T AND2T_38 (.a(net_r[48]), .b(net_r[329]), .clk(net_r[551]), .q(net_w[49]));
LSmitll_OR2T_v2p1_optimized OR2T_39 (.a(net_r[47]), .b(net_r[49]), .clk(net_r[557]), .q(net_w[50]));
LSmitll_XORT_v2p1_optimized XOR2T_40 (.a(net_r[46]), .b(net_r[330]), .clk(net_r[560]), .q(net_w[247]));
LSmitll_AND2T AND2T_41 (.a(net_r[277]), .b(net_r[308]), .clk(net_r[529]), .q(net_w[183]));
LSmitll_OR2T_v2p1_optimized OR2T_42 (.a(net_r[278]), .b(net_r[309]), .clk(net_r[528]), .q(net_w[52]));
LSmitll_AND2T AND2T_43 (.a(net_r[52]), .b(net_r[331]), .clk(net_r[562]), .q(net_w[53]));
LSmitll_OR2T_v2p1_optimized OR2T_44 (.a(net_r[51]), .b(net_r[53]), .clk(net_r[561]), .q(net_w[62]));
LSmitll_DFFT_v2p1_optimized DFF_71 (.a(net_r[63]), .clk(net_r[337]), .q(net_w[2]));
LSmitll_DFFT_v2p1_optimized DFF_72 (.a(net_r[64]), .clk(net_r[334]), .q(net_w[63]));
LSmitll_DFFT_v2p1_optimized DFF_73 (.a(net_r[65]), .clk(net_r[371]), .q(net_w[3]));
LSmitll_DFFT_v2p1_optimized DFF_74 (.a(net_r[66]), .clk(net_r[368]), .q(net_w[65]));
LSmitll_DFFT_v2p1_optimized DFF_75 (.a(net_r[67]), .clk(net_r[339]), .q(net_w[66]));
LSmitll_DFFT_v2p1_optimized DFF_76 (.a(net_r[68]), .clk(net_r[336]), .q(net_w[67]));
LSmitll_DFFT_v2p1_optimized DFF_77 (.a(net_r[69]), .clk(net_r[399]), .q(net_w[4]));
LSmitll_DFFT_v2p1_optimized DFF_78 (.a(net_r[70]), .clk(net_r[400]), .q(net_w[69]));
LSmitll_DFFT_v2p1_optimized DFF_79 (.a(net_r[71]), .clk(net_r[373]), .q(net_w[70]));
LSmitll_DFFT_v2p1_optimized DFF_80 (.a(net_r[72]), .clk(net_r[370]), .q(net_w[71]));
LSmitll_DFFT_v2p1_optimized DFF_81 (.a(net_r[73]), .clk(net_r[341]), .q(net_w[72]));
LSmitll_DFFT_v2p1_optimized DFF_82 (.a(net_r[74]), .clk(net_r[338]), .q(net_w[73]));
LSmitll_DFFT_v2p1_optimized DFF_83 (.a(net_r[75]), .clk(net_r[426]), .q(net_w[5]));
LSmitll_DFFT_v2p1_optimized DFF_84 (.a(net_r[76]), .clk(net_r[427]), .q(net_w[75]));
LSmitll_DFFT_v2p1_optimized DFF_85 (.a(net_r[77]), .clk(net_r[401]), .q(net_w[76]));
LSmitll_DFFT_v2p1_optimized DFF_86 (.a(net_r[78]), .clk(net_r[402]), .q(net_w[77]));
LSmitll_DFFT_v2p1_optimized DFF_87 (.a(net_r[79]), .clk(net_r[375]), .q(net_w[78]));
LSmitll_DFFT_v2p1_optimized DFF_88 (.a(net_r[80]), .clk(net_r[372]), .q(net_w[79]));
LSmitll_DFFT_v2p1_optimized DFF_89 (.a(net_r[81]), .clk(net_r[343]), .q(net_w[80]));
LSmitll_DFFT_v2p1_optimized DFF_90 (.a(net_r[82]), .clk(net_r[340]), .q(net_w[81]));
LSmitll_DFFT_v2p1_optimized DFF_91 (.a(net_r[83]), .clk(net_r[453]), .q(net_w[6]));
LSmitll_DFFT_v2p1_optimized DFF_92 (.a(net_r[84]), .clk(net_r[452]), .q(net_w[83]));
LSmitll_DFFT_v2p1_optimized DFF_93 (.a(net_r[85]), .clk(net_r[428]), .q(net_w[84]));
LSmitll_DFFT_v2p1_optimized DFF_94 (.a(net_r[86]), .clk(net_r[429]), .q(net_w[85]));
LSmitll_DFFT_v2p1_optimized DFF_95 (.a(net_r[87]), .clk(net_r[403]), .q(net_w[86]));
LSmitll_DFFT_v2p1_optimized DFF_96 (.a(net_r[88]), .clk(net_r[404]), .q(net_w[87]));
LSmitll_DFFT_v2p1_optimized DFF_97 (.a(net_r[89]), .clk(net_r[377]), .q(net_w[88]));
LSmitll_DFFT_v2p1_optimized DFF_98 (.a(net_r[90]), .clk(net_r[374]), .q(net_w[89]));
LSmitll_DFFT_v2p1_optimized DFF_99 (.a(net_r[91]), .clk(net_r[345]), .q(net_w[90]));
LSmitll_DFFT_v2p1_optimized DFF_100 (.a(net_r[92]), .clk(net_r[342]), .q(net_w[91]));
LSmitll_DFFT_v2p1_optimized DFF_101 (.a(net_r[93]), .clk(net_r[475]), .q(net_w[7]));
LSmitll_DFFT_v2p1_optimized DFF_102 (.a(net_r[94]), .clk(net_r[476]), .q(net_w[93]));
LSmitll_DFFT_v2p1_optimized DFF_103 (.a(net_r[95]), .clk(net_r[455]), .q(net_w[94]));
LSmitll_DFFT_v2p1_optimized DFF_104 (.a(net_r[96]), .clk(net_r[454]), .q(net_w[95]));
LSmitll_DFFT_v2p1_optimized DFF_105 (.a(net_r[97]), .clk(net_r[430]), .q(net_w[96]));
LSmitll_DFFT_v2p1_optimized DFF_106 (.a(net_r[98]), .clk(net_r[431]), .q(net_w[97]));
LSmitll_DFFT_v2p1_optimized DFF_107 (.a(net_r[99]), .clk(net_r[405]), .q(net_w[98]));
LSmitll_DFFT_v2p1_optimized DFF_108 (.a(net_r[100]), .clk(net_r[406]), .q(net_w[99]));
LSmitll_DFFT_v2p1_optimized DFF_109 (.a(net_r[101]), .clk(net_r[379]), .q(net_w[100]));
LSmitll_DFFT_v2p1_optimized DFF_110 (.a(net_r[102]), .clk(net_r[376]), .q(net_w[101]));
LSmitll_DFFT_v2p1_optimized DFF_111 (.a(net_r[103]), .clk(net_r[347]), .q(net_w[102]));
LSmitll_DFFT_v2p1_optimized DFF_112 (.a(net_r[104]), .clk(net_r[344]), .q(net_w[103]));
LSmitll_DFFT_v2p1_optimized DFF_113 (.a(net_r[105]), .clk(net_r[497]), .q(net_w[8]));
LSmitll_DFFT_v2p1_optimized DFF_114 (.a(net_r[106]), .clk(net_r[498]), .q(net_w[105]));
LSmitll_DFFT_v2p1_optimized DFF_115 (.a(net_r[107]), .clk(net_r[477]), .q(net_w[106]));
LSmitll_DFFT_v2p1_optimized DFF_116 (.a(net_r[108]), .clk(net_r[478]), .q(net_w[107]));
LSmitll_DFFT_v2p1_optimized DFF_117 (.a(net_r[109]), .clk(net_r[457]), .q(net_w[108]));
LSmitll_DFFT_v2p1_optimized DFF_118 (.a(net_r[110]), .clk(net_r[456]), .q(net_w[109]));
LSmitll_DFFT_v2p1_optimized DFF_119 (.a(net_r[111]), .clk(net_r[432]), .q(net_w[110]));
LSmitll_DFFT_v2p1_optimized DFF_120 (.a(net_r[112]), .clk(net_r[433]), .q(net_w[111]));
LSmitll_DFFT_v2p1_optimized DFF_121 (.a(net_r[113]), .clk(net_r[407]), .q(net_w[112]));
LSmitll_DFFT_v2p1_optimized DFF_122 (.a(net_r[114]), .clk(net_r[408]), .q(net_w[113]));
LSmitll_DFFT_v2p1_optimized DFF_123 (.a(net_r[115]), .clk(net_r[380]), .q(net_w[114]));
LSmitll_DFFT_v2p1_optimized DFF_124 (.a(net_r[116]), .clk(net_r[378]), .q(net_w[115]));
LSmitll_DFFT_v2p1_optimized DFF_125 (.a(net_r[117]), .clk(net_r[348]), .q(net_w[116]));
LSmitll_DFFT_v2p1_optimized DFF_126 (.a(net_r[118]), .clk(net_r[346]), .q(net_w[117]));
LSmitll_DFFT_v2p1_optimized DFF_127 (.a(net_r[119]), .clk(net_r[350]), .q(net_w[10]));
LSmitll_DFFT_v2p1_optimized DFF_128 (.a(net_r[120]), .clk(net_r[349]), .q(net_w[119]));
LSmitll_DFFT_v2p1_optimized DFF_129 (.a(net_r[121]), .clk(net_r[382]), .q(net_w[11]));
LSmitll_DFFT_v2p1_optimized DFF_130 (.a(net_r[122]), .clk(net_r[381]), .q(net_w[121]));
LSmitll_DFFT_v2p1_optimized DFF_131 (.a(net_r[123]), .clk(net_r[352]), .q(net_w[122]));
LSmitll_DFFT_v2p1_optimized DFF_132 (.a(net_r[124]), .clk(net_r[351]), .q(net_w[123]));
LSmitll_DFFT_v2p1_optimized DFF_133 (.a(net_r[125]), .clk(net_r[409]), .q(net_w[12]));
LSmitll_DFFT_v2p1_optimized DFF_134 (.a(net_r[126]), .clk(net_r[411]), .q(net_w[125]));
LSmitll_DFFT_v2p1_optimized DFF_135 (.a(net_r[127]), .clk(net_r[384]), .q(net_w[126]));
LSmitll_DFFT_v2p1_optimized DFF_136 (.a(net_r[128]), .clk(net_r[383]), .q(net_w[127]));
LSmitll_DFFT_v2p1_optimized DFF_137 (.a(net_r[129]), .clk(net_r[354]), .q(net_w[128]));
LSmitll_DFFT_v2p1_optimized DFF_138 (.a(net_r[130]), .clk(net_r[353]), .q(net_w[129]));
LSmitll_DFFT_v2p1_optimized DFF_139 (.a(net_r[131]), .clk(net_r[435]), .q(net_w[13]));
LSmitll_DFFT_v2p1_optimized DFF_140 (.a(net_r[132]), .clk(net_r[434]), .q(net_w[131]));
LSmitll_DFFT_v2p1_optimized DFF_141 (.a(net_r[133]), .clk(net_r[410]), .q(net_w[132]));
LSmitll_DFFT_v2p1_optimized DFF_142 (.a(net_r[134]), .clk(net_r[413]), .q(net_w[133]));
LSmitll_DFFT_v2p1_optimized DFF_143 (.a(net_r[135]), .clk(net_r[386]), .q(net_w[134]));
LSmitll_DFFT_v2p1_optimized DFF_144 (.a(net_r[136]), .clk(net_r[385]), .q(net_w[135]));
LSmitll_DFFT_v2p1_optimized DFF_145 (.a(net_r[137]), .clk(net_r[356]), .q(net_w[136]));
LSmitll_DFFT_v2p1_optimized DFF_146 (.a(net_r[138]), .clk(net_r[355]), .q(net_w[137]));
LSmitll_DFFT_v2p1_optimized DFF_147 (.a(net_r[139]), .clk(net_r[460]), .q(net_w[14]));
LSmitll_DFFT_v2p1_optimized DFF_148 (.a(net_r[140]), .clk(net_r[458]), .q(net_w[139]));
LSmitll_DFFT_v2p1_optimized DFF_149 (.a(net_r[141]), .clk(net_r[437]), .q(net_w[140]));
LSmitll_DFFT_v2p1_optimized DFF_150 (.a(net_r[142]), .clk(net_r[436]), .q(net_w[141]));
LSmitll_DFFT_v2p1_optimized DFF_151 (.a(net_r[143]), .clk(net_r[412]), .q(net_w[142]));
LSmitll_DFFT_v2p1_optimized DFF_152 (.a(net_r[144]), .clk(net_r[415]), .q(net_w[143]));
LSmitll_DFFT_v2p1_optimized DFF_153 (.a(net_r[145]), .clk(net_r[388]), .q(net_w[144]));
LSmitll_DFFT_v2p1_optimized DFF_154 (.a(net_r[146]), .clk(net_r[387]), .q(net_w[145]));
LSmitll_DFFT_v2p1_optimized DFF_155 (.a(net_r[147]), .clk(net_r[358]), .q(net_w[146]));
LSmitll_DFFT_v2p1_optimized DFF_156 (.a(net_r[148]), .clk(net_r[357]), .q(net_w[147]));
LSmitll_DFFT_v2p1_optimized DFF_157 (.a(net_r[149]), .clk(net_r[480]), .q(net_w[15]));
LSmitll_DFFT_v2p1_optimized DFF_158 (.a(net_r[150]), .clk(net_r[479]), .q(net_w[149]));
LSmitll_DFFT_v2p1_optimized DFF_159 (.a(net_r[151]), .clk(net_r[462]), .q(net_w[150]));
LSmitll_DFFT_v2p1_optimized DFF_160 (.a(net_r[152]), .clk(net_r[459]), .q(net_w[151]));
LSmitll_DFFT_v2p1_optimized DFF_161 (.a(net_r[153]), .clk(net_r[439]), .q(net_w[152]));
LSmitll_DFFT_v2p1_optimized DFF_162 (.a(net_r[154]), .clk(net_r[438]), .q(net_w[153]));
LSmitll_DFFT_v2p1_optimized DFF_163 (.a(net_r[155]), .clk(net_r[414]), .q(net_w[154]));
LSmitll_DFFT_v2p1_optimized DFF_164 (.a(net_r[156]), .clk(net_r[417]), .q(net_w[155]));
LSmitll_DFFT_v2p1_optimized DFF_165 (.a(net_r[157]), .clk(net_r[390]), .q(net_w[156]));
LSmitll_DFFT_v2p1_optimized DFF_166 (.a(net_r[158]), .clk(net_r[389]), .q(net_w[157]));
LSmitll_DFFT_v2p1_optimized DFF_167 (.a(net_r[159]), .clk(net_r[360]), .q(net_w[158]));
LSmitll_DFFT_v2p1_optimized DFF_168 (.a(net_r[160]), .clk(net_r[359]), .q(net_w[159]));
LSmitll_DFFT_v2p1_optimized DFF_169 (.a(net_r[161]), .clk(net_r[500]), .q(net_w[16]));
LSmitll_DFFT_v2p1_optimized DFF_170 (.a(net_r[162]), .clk(net_r[499]), .q(net_w[161]));
LSmitll_DFFT_v2p1_optimized DFF_171 (.a(net_r[163]), .clk(net_r[482]), .q(net_w[162]));
LSmitll_DFFT_v2p1_optimized DFF_172 (.a(net_r[164]), .clk(net_r[481]), .q(net_w[163]));
LSmitll_DFFT_v2p1_optimized DFF_173 (.a(net_r[165]), .clk(net_r[463]), .q(net_w[164]));
LSmitll_DFFT_v2p1_optimized DFF_174 (.a(net_r[166]), .clk(net_r[461]), .q(net_w[165]));
LSmitll_DFFT_v2p1_optimized DFF_175 (.a(net_r[167]), .clk(net_r[441]), .q(net_w[166]));
LSmitll_DFFT_v2p1_optimized DFF_176 (.a(net_r[168]), .clk(net_r[440]), .q(net_w[167]));
LSmitll_DFFT_v2p1_optimized DFF_177 (.a(net_r[169]), .clk(net_r[416]), .q(net_w[168]));
LSmitll_DFFT_v2p1_optimized DFF_178 (.a(net_r[170]), .clk(net_r[418]), .q(net_w[169]));
LSmitll_DFFT_v2p1_optimized DFF_179 (.a(net_r[171]), .clk(net_r[392]), .q(net_w[170]));
LSmitll_DFFT_v2p1_optimized DFF_180 (.a(net_r[172]), .clk(net_r[391]), .q(net_w[171]));
LSmitll_DFFT_v2p1_optimized DFF_181 (.a(net_r[173]), .clk(net_r[362]), .q(net_w[172]));
LSmitll_DFFT_v2p1_optimized DFF_182 (.a(net_r[174]), .clk(net_r[361]), .q(net_w[173]));
LSmitll_DFFT_v2p1_optimized DFF_183 (.a(net_r[175]), .clk(net_r[363]), .q(net_w[17]));
LSmitll_DFFT_v2p1_optimized DFF_184 (.a(net_r[176]), .clk(net_r[365]), .q(net_w[19]));
LSmitll_DFFT_v2p1_optimized DFF_185 (.a(net_r[177]), .clk(net_r[397]), .q(net_w[24]));
LSmitll_DFFT_v2p1_optimized DFF_186 (.a(net_r[178]), .clk(net_r[425]), .q(net_w[27]));
LSmitll_DFFT_v2p1_optimized DFF_187 (.a(net_r[179]), .clk(net_r[450]), .q(net_w[32]));
LSmitll_DFFT_v2p1_optimized DFF_188 (.a(net_r[180]), .clk(net_r[472]), .q(net_w[37]));
LSmitll_DFFT_v2p1_optimized DFF_189 (.a(net_r[181]), .clk(net_r[494]), .q(net_w[42]));
LSmitll_DFFT_v2p1_optimized DFF_190 (.a(net_r[182]), .clk(net_r[513]), .q(net_w[47]));
LSmitll_DFFT_v2p1_optimized DFF_191 (.a(net_r[183]), .clk(net_r[527]), .q(net_w[51]));
LSmitll_DFFT_v2p1_optimized DFF_192 (.a(net_r[184]), .clk(net_r[530]), .q(net_w[54]));
LSmitll_DFFT_v2p1_optimized DFF_193 (.a(net_r[185]), .clk(net_r[516]), .q(net_w[184]));
LSmitll_DFFT_v2p1_optimized DFF_194 (.a(net_r[186]), .clk(net_r[515]), .q(net_w[185]));
LSmitll_DFFT_v2p1_optimized DFF_195 (.a(net_r[187]), .clk(net_r[502]), .q(net_w[186]));
LSmitll_DFFT_v2p1_optimized DFF_196 (.a(net_r[188]), .clk(net_r[501]), .q(net_w[187]));
LSmitll_DFFT_v2p1_optimized DFF_197 (.a(net_r[189]), .clk(net_r[484]), .q(net_w[188]));
LSmitll_DFFT_v2p1_optimized DFF_198 (.a(net_r[190]), .clk(net_r[483]), .q(net_w[189]));
LSmitll_DFFT_v2p1_optimized DFF_199 (.a(net_r[191]), .clk(net_r[465]), .q(net_w[190]));
LSmitll_DFFT_v2p1_optimized DFF_200 (.a(net_r[192]), .clk(net_r[464]), .q(net_w[191]));
LSmitll_DFFT_v2p1_optimized DFF_201 (.a(net_r[193]), .clk(net_r[443]), .q(net_w[192]));
LSmitll_DFFT_v2p1_optimized DFF_202 (.a(net_r[194]), .clk(net_r[442]), .q(net_w[193]));
LSmitll_DFFT_v2p1_optimized DFF_203 (.a(net_r[195]), .clk(net_r[420]), .q(net_w[194]));
LSmitll_DFFT_v2p1_optimized DFF_204 (.a(net_r[196]), .clk(net_r[419]), .q(net_w[195]));
LSmitll_DFFT_v2p1_optimized DFF_205 (.a(net_r[197]), .clk(net_r[394]), .q(net_w[196]));
LSmitll_DFFT_v2p1_optimized DFF_206 (.a(net_r[198]), .clk(net_r[393]), .q(net_w[197]));
LSmitll_DFFT_v2p1_optimized DFF_207 (.a(net_r[199]), .clk(net_r[531]), .q(net_w[55]));
LSmitll_DFFT_v2p1_optimized DFF_208 (.a(net_r[200]), .clk(net_r[532]), .q(net_w[199]));
LSmitll_DFFT_v2p1_optimized DFF_209 (.a(net_r[201]), .clk(net_r[518]), .q(net_w[200]));
LSmitll_DFFT_v2p1_optimized DFF_210 (.a(net_r[202]), .clk(net_r[517]), .q(net_w[201]));
LSmitll_DFFT_v2p1_optimized DFF_211 (.a(net_r[203]), .clk(net_r[504]), .q(net_w[202]));
LSmitll_DFFT_v2p1_optimized DFF_212 (.a(net_r[204]), .clk(net_r[503]), .q(net_w[203]));
LSmitll_DFFT_v2p1_optimized DFF_213 (.a(net_r[205]), .clk(net_r[486]), .q(net_w[204]));
LSmitll_DFFT_v2p1_optimized DFF_214 (.a(net_r[206]), .clk(net_r[485]), .q(net_w[205]));
LSmitll_DFFT_v2p1_optimized DFF_215 (.a(net_r[207]), .clk(net_r[467]), .q(net_w[206]));
LSmitll_DFFT_v2p1_optimized DFF_216 (.a(net_r[208]), .clk(net_r[466]), .q(net_w[207]));
LSmitll_DFFT_v2p1_optimized DFF_217 (.a(net_r[209]), .clk(net_r[445]), .q(net_w[208]));
LSmitll_DFFT_v2p1_optimized DFF_218 (.a(net_r[210]), .clk(net_r[444]), .q(net_w[209]));
LSmitll_DFFT_v2p1_optimized DFF_219 (.a(net_r[211]), .clk(net_r[422]), .q(net_w[210]));
LSmitll_DFFT_v2p1_optimized DFF_220 (.a(net_r[212]), .clk(net_r[543]), .q(net_w[56]));
LSmitll_DFFT_v2p1_optimized DFF_221 (.a(net_r[213]), .clk(net_r[533]), .q(net_w[212]));
LSmitll_DFFT_v2p1_optimized DFF_222 (.a(net_r[214]), .clk(net_r[534]), .q(net_w[213]));
LSmitll_DFFT_v2p1_optimized DFF_223 (.a(net_r[215]), .clk(net_r[520]), .q(net_w[214]));
LSmitll_DFFT_v2p1_optimized DFF_224 (.a(net_r[216]), .clk(net_r[519]), .q(net_w[215]));
LSmitll_DFFT_v2p1_optimized DFF_225 (.a(net_r[217]), .clk(net_r[506]), .q(net_w[216]));
LSmitll_DFFT_v2p1_optimized DFF_226 (.a(net_r[218]), .clk(net_r[505]), .q(net_w[217]));
LSmitll_DFFT_v2p1_optimized DFF_227 (.a(net_r[219]), .clk(net_r[488]), .q(net_w[218]));
LSmitll_DFFT_v2p1_optimized DFF_228 (.a(net_r[220]), .clk(net_r[487]), .q(net_w[219]));
LSmitll_DFFT_v2p1_optimized DFF_229 (.a(net_r[221]), .clk(net_r[469]), .q(net_w[220]));
LSmitll_DFFT_v2p1_optimized DFF_230 (.a(net_r[222]), .clk(net_r[468]), .q(net_w[221]));
LSmitll_DFFT_v2p1_optimized DFF_231 (.a(net_r[223]), .clk(net_r[544]), .q(net_w[57]));
LSmitll_DFFT_v2p1_optimized DFF_232 (.a(net_r[224]), .clk(net_r[545]), .q(net_w[223]));
LSmitll_DFFT_v2p1_optimized DFF_233 (.a(net_r[225]), .clk(net_r[535]), .q(net_w[224]));
LSmitll_DFFT_v2p1_optimized DFF_234 (.a(net_r[226]), .clk(net_r[536]), .q(net_w[225]));
LSmitll_DFFT_v2p1_optimized DFF_235 (.a(net_r[227]), .clk(net_r[522]), .q(net_w[226]));
LSmitll_DFFT_v2p1_optimized DFF_236 (.a(net_r[228]), .clk(net_r[521]), .q(net_w[227]));
LSmitll_DFFT_v2p1_optimized DFF_237 (.a(net_r[229]), .clk(net_r[508]), .q(net_w[228]));
LSmitll_DFFT_v2p1_optimized DFF_238 (.a(net_r[230]), .clk(net_r[507]), .q(net_w[229]));
LSmitll_DFFT_v2p1_optimized DFF_239 (.a(net_r[231]), .clk(net_r[490]), .q(net_w[230]));
LSmitll_DFFT_v2p1_optimized DFF_240 (.a(net_r[232]), .clk(net_r[552]), .q(net_w[58]));
LSmitll_DFFT_v2p1_optimized DFF_241 (.a(net_r[233]), .clk(net_r[546]), .q(net_w[232]));
LSmitll_DFFT_v2p1_optimized DFF_242 (.a(net_r[234]), .clk(net_r[547]), .q(net_w[233]));
LSmitll_DFFT_v2p1_optimized DFF_243 (.a(net_r[235]), .clk(net_r[537]), .q(net_w[234]));
LSmitll_DFFT_v2p1_optimized DFF_244 (.a(net_r[236]), .clk(net_r[538]), .q(net_w[235]));
LSmitll_DFFT_v2p1_optimized DFF_245 (.a(net_r[237]), .clk(net_r[524]), .q(net_w[236]));
LSmitll_DFFT_v2p1_optimized DFF_246 (.a(net_r[238]), .clk(net_r[523]), .q(net_w[237]));
LSmitll_DFFT_v2p1_optimized DFF_247 (.a(net_r[239]), .clk(net_r[553]), .q(net_w[59]));
LSmitll_DFFT_v2p1_optimized DFF_248 (.a(net_r[240]), .clk(net_r[554]), .q(net_w[239]));
LSmitll_DFFT_v2p1_optimized DFF_249 (.a(net_r[241]), .clk(net_r[548]), .q(net_w[240]));
LSmitll_DFFT_v2p1_optimized DFF_250 (.a(net_r[242]), .clk(net_r[549]), .q(net_w[241]));
LSmitll_DFFT_v2p1_optimized DFF_251 (.a(net_r[243]), .clk(net_r[539]), .q(net_w[242]));
LSmitll_DFFT_v2p1_optimized DFF_252 (.a(net_r[244]), .clk(net_r[558]), .q(net_w[60]));
LSmitll_DFFT_v2p1_optimized DFF_253 (.a(net_r[245]), .clk(net_r[555]), .q(net_w[244]));
LSmitll_DFFT_v2p1_optimized DFF_254 (.a(net_r[246]), .clk(net_r[556]), .q(net_w[245]));
LSmitll_DFFT_v2p1_optimized DFF_255 (.a(net_r[247]), .clk(net_r[559]), .q(net_w[61]));
LSmitll_SPLITT_v2p1_optimized SPLIT_256 (.a(net_r[1]), .q(net_w[248]), .m(net_w[249]));
LSmitll_SPLITT_v2p1_optimized SPLIT_257 (.a(net_r[2]), .q(net_w[250]), .m(net_w[251]));
LSmitll_SPLITT_v2p1_optimized SPLIT_258 (.a(net_r[3]), .q(net_w[252]), .m(net_w[253]));
LSmitll_SPLITT_v2p1_optimized SPLIT_259 (.a(net_r[4]), .q(net_w[254]), .m(net_w[255]));
LSmitll_SPLITT_v2p1_optimized SPLIT_260 (.a(net_r[254]), .q(net_w[256]), .m(net_w[258]));
LSmitll_SPLITT_v2p1_optimized SPLIT_261 (.a(net_r[255]), .q(net_w[257]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_262 (.a(net_r[5]), .q(net_w[259]), .m(net_w[260]));
LSmitll_SPLITT_v2p1_optimized SPLIT_263 (.a(net_r[259]), .q(net_w[261]), .m(net_w[263]));
LSmitll_SPLITT_v2p1_optimized SPLIT_264 (.a(net_r[260]), .q(net_w[262]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_265 (.a(net_r[6]), .q(net_w[264]), .m(net_w[265]));
LSmitll_SPLITT_v2p1_optimized SPLIT_266 (.a(net_r[264]), .q(net_w[266]), .m(net_w[268]));
LSmitll_SPLITT_v2p1_optimized SPLIT_267 (.a(net_r[265]), .q(net_w[267]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_268 (.a(net_r[7]), .q(net_w[269]), .m(net_w[270]));
LSmitll_SPLITT_v2p1_optimized SPLIT_269 (.a(net_r[269]), .q(net_w[271]), .m(net_w[273]));
LSmitll_SPLITT_v2p1_optimized SPLIT_270 (.a(net_r[270]), .q(net_w[272]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_271 (.a(net_r[8]), .q(net_w[274]), .m(net_w[275]));
LSmitll_SPLITT_v2p1_optimized SPLIT_272 (.a(net_r[274]), .q(net_w[276]), .m(net_w[278]));
LSmitll_SPLITT_v2p1_optimized SPLIT_273 (.a(net_r[275]), .q(net_w[277]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_274 (.a(net_r[9]), .q(net_w[279]), .m(net_w[280]));
LSmitll_SPLITT_v2p1_optimized SPLIT_275 (.a(net_r[10]), .q(net_w[281]), .m(net_w[282]));
LSmitll_SPLITT_v2p1_optimized SPLIT_276 (.a(net_r[11]), .q(net_w[283]), .m(net_w[284]));
LSmitll_SPLITT_v2p1_optimized SPLIT_277 (.a(net_r[12]), .q(net_w[285]), .m(net_w[286]));
LSmitll_SPLITT_v2p1_optimized SPLIT_278 (.a(net_r[285]), .q(net_w[287]), .m(net_w[289]));
LSmitll_SPLITT_v2p1_optimized SPLIT_279 (.a(net_r[286]), .q(net_w[288]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_280 (.a(net_r[13]), .q(net_w[290]), .m(net_w[291]));
LSmitll_SPLITT_v2p1_optimized SPLIT_281 (.a(net_r[290]), .q(net_w[292]), .m(net_w[294]));
LSmitll_SPLITT_v2p1_optimized SPLIT_282 (.a(net_r[291]), .q(net_w[293]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_283 (.a(net_r[14]), .q(net_w[295]), .m(net_w[296]));
LSmitll_SPLITT_v2p1_optimized SPLIT_284 (.a(net_r[295]), .q(net_w[297]), .m(net_w[299]));
LSmitll_SPLITT_v2p1_optimized SPLIT_285 (.a(net_r[296]), .q(net_w[298]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_286 (.a(net_r[15]), .q(net_w[300]), .m(net_w[301]));
LSmitll_SPLITT_v2p1_optimized SPLIT_287 (.a(net_r[300]), .q(net_w[302]), .m(net_w[304]));
LSmitll_SPLITT_v2p1_optimized SPLIT_288 (.a(net_r[301]), .q(net_w[303]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_289 (.a(net_r[16]), .q(net_w[305]), .m(net_w[306]));
LSmitll_SPLITT_v2p1_optimized SPLIT_290 (.a(net_r[305]), .q(net_w[307]), .m(net_w[309]));
LSmitll_SPLITT_v2p1_optimized SPLIT_291 (.a(net_r[306]), .q(net_w[308]), .m());
LSmitll_SPLITT_v2p1_optimized SPLIT_292 (.a(net_r[17]), .q(net_w[310]), .m(net_w[311]));
LSmitll_SPLITT_v2p1_optimized SPLIT_293 (.a(net_r[18]), .q(net_w[312]), .m(net_w[313]));
LSmitll_SPLITT_v2p1_optimized SPLIT_294 (.a(net_r[21]), .q(net_w[314]), .m(net_w[315]));
LSmitll_SPLITT_v2p1_optimized SPLIT_295 (.a(net_r[22]), .q(net_w[316]), .m(net_w[317]));
LSmitll_SPLITT_v2p1_optimized SPLIT_296 (.a(net_r[23]), .q(net_w[318]), .m(net_w[319]));
LSmitll_SPLITT_v2p1_optimized SPLIT_297 (.a(net_r[26]), .q(net_w[320]), .m(net_w[321]));
LSmitll_SPLITT_v2p1_optimized SPLIT_298 (.a(net_r[29]), .q(net_w[322]), .m(net_w[323]));
LSmitll_SPLITT_v2p1_optimized SPLIT_299 (.a(net_r[35]), .q(net_w[324]), .m(net_w[325]));
LSmitll_SPLITT_v2p1_optimized SPLIT_300 (.a(net_r[40]), .q(net_w[326]), .m(net_w[327]));
LSmitll_SPLITT_v2p1_optimized SPLIT_301 (.a(net_r[45]), .q(net_w[328]), .m(net_w[329]));
LSmitll_SPLITT_v2p1_optimized SPLIT_302 (.a(net_r[50]), .q(net_w[330]), .m(net_w[331]));
LSmitll_SPLITT_v2p1_optimized SC_304 (.a(net_r[563]), .q(net_w[333]), .m(net_w[334]));
LSmitll_SPLITT_v2p1_optimized SC_305 (.a(net_r[564]), .q(net_w[335]), .m(net_w[336]));
LSmitll_SPLITT_v2p1_optimized SC_306 (.a(net_r[565]), .q(net_w[337]), .m(net_w[338]));
LSmitll_SPLITT_v2p1_optimized SC_307 (.a(net_r[566]), .q(net_w[339]), .m(net_w[340]));
LSmitll_SPLITT_v2p1_optimized SC_308 (.a(net_r[567]), .q(net_w[341]), .m(net_w[342]));
LSmitll_SPLITT_v2p1_optimized SC_309 (.a(net_r[568]), .q(net_w[343]), .m(net_w[344]));
LSmitll_SPLITT_v2p1_optimized SC_310 (.a(net_r[569]), .q(net_w[345]), .m(net_w[346]));
LSmitll_SPLITT_v2p1_optimized SC_311 (.a(net_r[570]), .q(net_w[347]), .m(net_w[348]));
LSmitll_SPLITT_v2p1_optimized SC_312 (.a(net_r[571]), .q(net_w[349]), .m(net_w[350]));
LSmitll_SPLITT_v2p1_optimized SC_313 (.a(net_r[572]), .q(net_w[351]), .m(net_w[352]));
LSmitll_SPLITT_v2p1_optimized SC_314 (.a(net_r[573]), .q(net_w[353]), .m(net_w[354]));
LSmitll_SPLITT_v2p1_optimized SC_315 (.a(net_r[574]), .q(net_w[355]), .m(net_w[356]));
LSmitll_SPLITT_v2p1_optimized SC_316 (.a(net_r[575]), .q(net_w[357]), .m(net_w[358]));
LSmitll_SPLITT_v2p1_optimized SC_317 (.a(net_r[576]), .q(net_w[359]), .m(net_w[360]));
LSmitll_SPLITT_v2p1_optimized SC_318 (.a(net_r[577]), .q(net_w[361]), .m(net_w[362]));
LSmitll_SPLITT_v2p1_optimized SC_319 (.a(net_r[578]), .q(net_w[363]), .m());
LSmitll_SPLITT_v2p1_optimized SC_320 (.a(net_r[593]), .q(net_w[364]), .m(net_w[365]));
LSmitll_SPLITT_v2p1_optimized SC_321 (.a(net_r[594]), .q(net_w[366]), .m(net_w[367]));
LSmitll_SPLITT_v2p1_optimized SC_322 (.a(net_r[595]), .q(net_w[368]), .m(net_w[369]));
LSmitll_SPLITT_v2p1_optimized SC_323 (.a(net_r[596]), .q(net_w[370]), .m(net_w[371]));
LSmitll_SPLITT_v2p1_optimized SC_324 (.a(net_r[597]), .q(net_w[372]), .m(net_w[373]));
LSmitll_SPLITT_v2p1_optimized SC_325 (.a(net_r[598]), .q(net_w[374]), .m(net_w[375]));
LSmitll_SPLITT_v2p1_optimized SC_326 (.a(net_r[599]), .q(net_w[376]), .m(net_w[377]));
LSmitll_SPLITT_v2p1_optimized SC_327 (.a(net_r[600]), .q(net_w[378]), .m(net_w[379]));
LSmitll_SPLITT_v2p1_optimized SC_328 (.a(net_r[601]), .q(net_w[380]), .m(net_w[381]));
LSmitll_SPLITT_v2p1_optimized SC_329 (.a(net_r[602]), .q(net_w[382]), .m(net_w[383]));
LSmitll_SPLITT_v2p1_optimized SC_330 (.a(net_r[603]), .q(net_w[384]), .m(net_w[385]));
LSmitll_SPLITT_v2p1_optimized SC_331 (.a(net_r[604]), .q(net_w[386]), .m(net_w[387]));
LSmitll_SPLITT_v2p1_optimized SC_332 (.a(net_r[605]), .q(net_w[388]), .m(net_w[389]));
LSmitll_SPLITT_v2p1_optimized SC_333 (.a(net_r[606]), .q(net_w[390]), .m(net_w[391]));
LSmitll_SPLITT_v2p1_optimized SC_334 (.a(net_r[607]), .q(net_w[392]), .m());
LSmitll_SPLITT_v2p1_optimized SC_335 (.a(net_r[622]), .q(net_w[393]), .m(net_w[394]));
LSmitll_SPLITT_v2p1_optimized SC_336 (.a(net_r[623]), .q(net_w[395]), .m(net_w[396]));
LSmitll_SPLITT_v2p1_optimized SC_337 (.a(net_r[624]), .q(net_w[397]), .m(net_w[398]));
LSmitll_SPLITT_v2p1_optimized SC_338 (.a(net_r[625]), .q(net_w[399]), .m(net_w[400]));
LSmitll_SPLITT_v2p1_optimized SC_339 (.a(net_r[626]), .q(net_w[401]), .m(net_w[402]));
LSmitll_SPLITT_v2p1_optimized SC_340 (.a(net_r[627]), .q(net_w[403]), .m(net_w[404]));
LSmitll_SPLITT_v2p1_optimized SC_341 (.a(net_r[628]), .q(net_w[405]), .m(net_w[406]));
LSmitll_SPLITT_v2p1_optimized SC_342 (.a(net_r[629]), .q(net_w[407]), .m(net_w[408]));
LSmitll_SPLITT_v2p1_optimized SC_343 (.a(net_r[630]), .q(net_w[409]), .m(net_w[410]));
LSmitll_SPLITT_v2p1_optimized SC_344 (.a(net_r[631]), .q(net_w[411]), .m(net_w[412]));
LSmitll_SPLITT_v2p1_optimized SC_345 (.a(net_r[632]), .q(net_w[413]), .m(net_w[414]));
LSmitll_SPLITT_v2p1_optimized SC_346 (.a(net_r[633]), .q(net_w[415]), .m(net_w[416]));
LSmitll_SPLITT_v2p1_optimized SC_347 (.a(net_r[634]), .q(net_w[417]), .m(net_w[418]));
LSmitll_SPLITT_v2p1_optimized SC_348 (.a(net_r[648]), .q(net_w[419]), .m(net_w[420]));
LSmitll_SPLITT_v2p1_optimized SC_349 (.a(net_r[649]), .q(net_w[421]), .m(net_w[422]));
LSmitll_SPLITT_v2p1_optimized SC_350 (.a(net_r[650]), .q(net_w[423]), .m(net_w[424]));
LSmitll_SPLITT_v2p1_optimized SC_351 (.a(net_r[651]), .q(net_w[425]), .m(net_w[426]));
LSmitll_SPLITT_v2p1_optimized SC_352 (.a(net_r[652]), .q(net_w[427]), .m(net_w[428]));
LSmitll_SPLITT_v2p1_optimized SC_353 (.a(net_r[653]), .q(net_w[429]), .m(net_w[430]));
LSmitll_SPLITT_v2p1_optimized SC_354 (.a(net_r[654]), .q(net_w[431]), .m(net_w[432]));
LSmitll_SPLITT_v2p1_optimized SC_355 (.a(net_r[655]), .q(net_w[433]), .m(net_w[434]));
LSmitll_SPLITT_v2p1_optimized SC_356 (.a(net_r[656]), .q(net_w[435]), .m(net_w[436]));
LSmitll_SPLITT_v2p1_optimized SC_357 (.a(net_r[657]), .q(net_w[437]), .m(net_w[438]));
LSmitll_SPLITT_v2p1_optimized SC_358 (.a(net_r[658]), .q(net_w[439]), .m(net_w[440]));
LSmitll_SPLITT_v2p1_optimized SC_359 (.a(net_r[659]), .q(net_w[441]), .m());
LSmitll_SPLITT_v2p1_optimized SC_360 (.a(net_r[671]), .q(net_w[442]), .m(net_w[443]));
LSmitll_SPLITT_v2p1_optimized SC_361 (.a(net_r[672]), .q(net_w[444]), .m(net_w[445]));
LSmitll_SPLITT_v2p1_optimized SC_362 (.a(net_r[673]), .q(net_w[446]), .m(net_w[447]));
LSmitll_SPLITT_v2p1_optimized SC_363 (.a(net_r[674]), .q(net_w[448]), .m(net_w[449]));
LSmitll_SPLITT_v2p1_optimized SC_364 (.a(net_r[675]), .q(net_w[450]), .m(net_w[451]));
LSmitll_SPLITT_v2p1_optimized SC_365 (.a(net_r[676]), .q(net_w[452]), .m(net_w[453]));
LSmitll_SPLITT_v2p1_optimized SC_366 (.a(net_r[677]), .q(net_w[454]), .m(net_w[455]));
LSmitll_SPLITT_v2p1_optimized SC_367 (.a(net_r[678]), .q(net_w[456]), .m(net_w[457]));
LSmitll_SPLITT_v2p1_optimized SC_368 (.a(net_r[679]), .q(net_w[458]), .m(net_w[459]));
LSmitll_SPLITT_v2p1_optimized SC_369 (.a(net_r[680]), .q(net_w[460]), .m(net_w[461]));
LSmitll_SPLITT_v2p1_optimized SC_370 (.a(net_r[681]), .q(net_w[462]), .m(net_w[463]));
LSmitll_SPLITT_v2p1_optimized SC_371 (.a(net_r[693]), .q(net_w[464]), .m(net_w[465]));
LSmitll_SPLITT_v2p1_optimized SC_372 (.a(net_r[694]), .q(net_w[466]), .m(net_w[467]));
LSmitll_SPLITT_v2p1_optimized SC_373 (.a(net_r[695]), .q(net_w[468]), .m(net_w[469]));
LSmitll_SPLITT_v2p1_optimized SC_374 (.a(net_r[696]), .q(net_w[470]), .m(net_w[471]));
LSmitll_SPLITT_v2p1_optimized SC_375 (.a(net_r[697]), .q(net_w[472]), .m(net_w[473]));
LSmitll_SPLITT_v2p1_optimized SC_376 (.a(net_r[698]), .q(net_w[474]), .m(net_w[475]));
LSmitll_SPLITT_v2p1_optimized SC_377 (.a(net_r[699]), .q(net_w[476]), .m(net_w[477]));
LSmitll_SPLITT_v2p1_optimized SC_378 (.a(net_r[700]), .q(net_w[478]), .m(net_w[479]));
LSmitll_SPLITT_v2p1_optimized SC_379 (.a(net_r[701]), .q(net_w[480]), .m(net_w[481]));
LSmitll_SPLITT_v2p1_optimized SC_380 (.a(net_r[702]), .q(net_w[482]), .m());
LSmitll_SPLITT_v2p1_optimized SC_381 (.a(net_r[713]), .q(net_w[483]), .m(net_w[484]));
LSmitll_SPLITT_v2p1_optimized SC_382 (.a(net_r[714]), .q(net_w[485]), .m(net_w[486]));
LSmitll_SPLITT_v2p1_optimized SC_383 (.a(net_r[715]), .q(net_w[487]), .m(net_w[488]));
LSmitll_SPLITT_v2p1_optimized SC_384 (.a(net_r[716]), .q(net_w[489]), .m(net_w[490]));
LSmitll_SPLITT_v2p1_optimized SC_385 (.a(net_r[717]), .q(net_w[491]), .m(net_w[492]));
LSmitll_SPLITT_v2p1_optimized SC_386 (.a(net_r[718]), .q(net_w[493]), .m(net_w[494]));
LSmitll_SPLITT_v2p1_optimized SC_387 (.a(net_r[719]), .q(net_w[495]), .m(net_w[496]));
LSmitll_SPLITT_v2p1_optimized SC_388 (.a(net_r[720]), .q(net_w[497]), .m(net_w[498]));
LSmitll_SPLITT_v2p1_optimized SC_389 (.a(net_r[721]), .q(net_w[499]), .m(net_w[500]));
LSmitll_SPLITT_v2p1_optimized SC_390 (.a(net_r[732]), .q(net_w[501]), .m(net_w[502]));
LSmitll_SPLITT_v2p1_optimized SC_391 (.a(net_r[733]), .q(net_w[503]), .m(net_w[504]));
LSmitll_SPLITT_v2p1_optimized SC_392 (.a(net_r[734]), .q(net_w[505]), .m(net_w[506]));
LSmitll_SPLITT_v2p1_optimized SC_393 (.a(net_r[735]), .q(net_w[507]), .m(net_w[508]));
LSmitll_SPLITT_v2p1_optimized SC_394 (.a(net_r[736]), .q(net_w[509]), .m(net_w[510]));
LSmitll_SPLITT_v2p1_optimized SC_395 (.a(net_r[737]), .q(net_w[511]), .m(net_w[512]));
LSmitll_SPLITT_v2p1_optimized SC_396 (.a(net_r[738]), .q(net_w[513]), .m(net_w[514]));
LSmitll_SPLITT_v2p1_optimized SC_397 (.a(net_r[746]), .q(net_w[515]), .m(net_w[516]));
LSmitll_SPLITT_v2p1_optimized SC_398 (.a(net_r[747]), .q(net_w[517]), .m(net_w[518]));
LSmitll_SPLITT_v2p1_optimized SC_399 (.a(net_r[748]), .q(net_w[519]), .m(net_w[520]));
LSmitll_SPLITT_v2p1_optimized SC_400 (.a(net_r[749]), .q(net_w[521]), .m(net_w[522]));
LSmitll_SPLITT_v2p1_optimized SC_401 (.a(net_r[750]), .q(net_w[523]), .m(net_w[524]));
LSmitll_SPLITT_v2p1_optimized SC_402 (.a(net_r[751]), .q(net_w[525]), .m(net_w[526]));
LSmitll_SPLITT_v2p1_optimized SC_403 (.a(net_r[752]), .q(net_w[527]), .m(net_w[528]));
LSmitll_SPLITT_v2p1_optimized SC_404 (.a(net_r[753]), .q(net_w[529]), .m());
LSmitll_SPLITT_v2p1_optimized SC_405 (.a(net_r[761]), .q(net_w[530]), .m(net_w[531]));
LSmitll_SPLITT_v2p1_optimized SC_406 (.a(net_r[762]), .q(net_w[532]), .m(net_w[533]));
LSmitll_SPLITT_v2p1_optimized SC_407 (.a(net_r[763]), .q(net_w[534]), .m(net_w[535]));
LSmitll_SPLITT_v2p1_optimized SC_408 (.a(net_r[764]), .q(net_w[536]), .m(net_w[537]));
LSmitll_SPLITT_v2p1_optimized SC_409 (.a(net_r[765]), .q(net_w[538]), .m(net_w[539]));
LSmitll_SPLITT_v2p1_optimized SC_410 (.a(net_r[766]), .q(net_w[540]), .m(net_w[541]));
LSmitll_SPLITT_v2p1_optimized SC_411 (.a(net_r[767]), .q(net_w[542]), .m());
LSmitll_SPLITT_v2p1_optimized SC_412 (.a(net_r[775]), .q(net_w[543]), .m(net_w[544]));
LSmitll_SPLITT_v2p1_optimized SC_413 (.a(net_r[776]), .q(net_w[545]), .m(net_w[546]));
LSmitll_SPLITT_v2p1_optimized SC_414 (.a(net_r[777]), .q(net_w[547]), .m(net_w[548]));
LSmitll_SPLITT_v2p1_optimized SC_415 (.a(net_r[778]), .q(net_w[549]), .m(net_w[550]));
LSmitll_SPLITT_v2p1_optimized SC_416 (.a(net_r[779]), .q(net_w[551]), .m());
LSmitll_SPLITT_v2p1_optimized SC_417 (.a(net_r[786]), .q(net_w[552]), .m(net_w[553]));
LSmitll_SPLITT_v2p1_optimized SC_418 (.a(net_r[787]), .q(net_w[554]), .m(net_w[555]));
LSmitll_SPLITT_v2p1_optimized SC_419 (.a(net_r[788]), .q(net_w[556]), .m(net_w[557]));
LSmitll_SPLITT_v2p1_optimized SC_420 (.a(net_r[793]), .q(net_w[558]), .m(net_w[559]));
LSmitll_SPLITT_v2p1_optimized SC_421 (.a(net_r[794]), .q(net_w[560]), .m(net_w[561]));
LSmitll_SPLITT_v2p1_optimized SC_422 (.a(net_r[795]), .q(net_w[562]), .m());
LSmitll_SPLITT_v2p1_optimized SC_423 (.a(net_r[579]), .q(net_w[563]), .m(net_w[564]));
LSmitll_SPLITT_v2p1_optimized SC_424 (.a(net_r[580]), .q(net_w[565]), .m(net_w[566]));
LSmitll_SPLITT_v2p1_optimized SC_425 (.a(net_r[581]), .q(net_w[567]), .m(net_w[568]));
LSmitll_SPLITT_v2p1_optimized SC_426 (.a(net_r[582]), .q(net_w[569]), .m(net_w[570]));
LSmitll_SPLITT_v2p1_optimized SC_427 (.a(net_r[583]), .q(net_w[571]), .m(net_w[572]));
LSmitll_SPLITT_v2p1_optimized SC_428 (.a(net_r[584]), .q(net_w[573]), .m(net_w[574]));
LSmitll_SPLITT_v2p1_optimized SC_429 (.a(net_r[585]), .q(net_w[575]), .m(net_w[576]));
LSmitll_SPLITT_v2p1_optimized SC_430 (.a(net_r[586]), .q(net_w[577]), .m(net_w[578]));
LSmitll_SPLITT_v2p1_optimized SC_431 (.a(net_r[587]), .q(net_w[579]), .m(net_w[580]));
LSmitll_SPLITT_v2p1_optimized SC_432 (.a(net_r[588]), .q(net_w[581]), .m(net_w[582]));
LSmitll_SPLITT_v2p1_optimized SC_433 (.a(net_r[589]), .q(net_w[583]), .m(net_w[584]));
LSmitll_SPLITT_v2p1_optimized SC_434 (.a(net_r[590]), .q(net_w[585]), .m(net_w[586]));
LSmitll_SPLITT_v2p1_optimized SC_435 (.a(net_r[591]), .q(net_w[587]), .m(net_w[588]));
LSmitll_SPLITT_v2p1_optimized SC_436 (.a(net_r[592]), .q(net_w[589]), .m(net_w[590]));
LSmitll_SPLITT_v2p1_optimized SC_437 (.a(net_r[814]), .q(net_w[591]), .m(net_w[592]));
LSmitll_SPLITT_v2p1_optimized SC_438 (.a(net_r[608]), .q(net_w[593]), .m(net_w[594]));
LSmitll_SPLITT_v2p1_optimized SC_439 (.a(net_r[609]), .q(net_w[595]), .m(net_w[596]));
LSmitll_SPLITT_v2p1_optimized SC_440 (.a(net_r[610]), .q(net_w[597]), .m(net_w[598]));
LSmitll_SPLITT_v2p1_optimized SC_441 (.a(net_r[611]), .q(net_w[599]), .m(net_w[600]));
LSmitll_SPLITT_v2p1_optimized SC_442 (.a(net_r[613]), .q(net_w[601]), .m(net_w[602]));
LSmitll_SPLITT_v2p1_optimized SC_443 (.a(net_r[614]), .q(net_w[603]), .m(net_w[604]));
LSmitll_SPLITT_v2p1_optimized SC_444 (.a(net_r[615]), .q(net_w[605]), .m(net_w[606]));
LSmitll_SPLITT_v2p1_optimized SC_445 (.a(net_r[612]), .q(net_w[607]), .m());
LSmitll_SPLITT_v2p1_optimized SC_446 (.a(net_r[616]), .q(net_w[608]), .m(net_w[609]));
LSmitll_SPLITT_v2p1_optimized SC_447 (.a(net_r[617]), .q(net_w[610]), .m(net_w[611]));
LSmitll_SPLITT_v2p1_optimized SC_448 (.a(net_r[618]), .q(net_w[612]), .m(net_w[613]));
LSmitll_SPLITT_v2p1_optimized SC_449 (.a(net_r[619]), .q(net_w[614]), .m(net_w[615]));
LSmitll_SPLITT_v2p1_optimized SC_450 (.a(net_r[620]), .q(net_w[616]), .m(net_w[617]));
LSmitll_SPLITT_v2p1_optimized SC_451 (.a(net_r[621]), .q(net_w[618]), .m(net_w[619]));
LSmitll_SPLITT_v2p1_optimized SC_452 (.a(net_r[815]), .q(net_w[620]), .m(net_w[621]));
LSmitll_SPLITT_v2p1_optimized SC_453 (.a(net_r[635]), .q(net_w[622]), .m(net_w[623]));
LSmitll_SPLITT_v2p1_optimized SC_454 (.a(net_r[636]), .q(net_w[624]), .m(net_w[625]));
LSmitll_SPLITT_v2p1_optimized SC_455 (.a(net_r[637]), .q(net_w[626]), .m(net_w[627]));
LSmitll_SPLITT_v2p1_optimized SC_456 (.a(net_r[638]), .q(net_w[628]), .m(net_w[629]));
LSmitll_SPLITT_v2p1_optimized SC_457 (.a(net_r[640]), .q(net_w[630]), .m(net_w[631]));
LSmitll_SPLITT_v2p1_optimized SC_458 (.a(net_r[641]), .q(net_w[632]), .m(net_w[633]));
LSmitll_SPLITT_v2p1_optimized SC_459 (.a(net_r[639]), .q(net_w[634]), .m());
LSmitll_SPLITT_v2p1_optimized SC_460 (.a(net_r[642]), .q(net_w[635]), .m(net_w[636]));
LSmitll_SPLITT_v2p1_optimized SC_461 (.a(net_r[643]), .q(net_w[637]), .m(net_w[638]));
LSmitll_SPLITT_v2p1_optimized SC_462 (.a(net_r[645]), .q(net_w[639]), .m(net_w[640]));
LSmitll_SPLITT_v2p1_optimized SC_463 (.a(net_r[644]), .q(net_w[641]), .m());
LSmitll_SPLITT_v2p1_optimized SC_464 (.a(net_r[646]), .q(net_w[642]), .m(net_w[643]));
LSmitll_SPLITT_v2p1_optimized SC_465 (.a(net_r[647]), .q(net_w[644]), .m(net_w[645]));
LSmitll_SPLITT_v2p1_optimized SC_466 (.a(net_r[816]), .q(net_w[646]), .m(net_w[647]));
LSmitll_SPLITT_v2p1_optimized SC_467 (.a(net_r[660]), .q(net_w[648]), .m(net_w[649]));
LSmitll_SPLITT_v2p1_optimized SC_468 (.a(net_r[661]), .q(net_w[650]), .m(net_w[651]));
LSmitll_SPLITT_v2p1_optimized SC_469 (.a(net_r[662]), .q(net_w[652]), .m(net_w[653]));
LSmitll_SPLITT_v2p1_optimized SC_470 (.a(net_r[663]), .q(net_w[654]), .m(net_w[655]));
LSmitll_SPLITT_v2p1_optimized SC_471 (.a(net_r[664]), .q(net_w[656]), .m(net_w[657]));
LSmitll_SPLITT_v2p1_optimized SC_472 (.a(net_r[665]), .q(net_w[658]), .m(net_w[659]));
LSmitll_SPLITT_v2p1_optimized SC_473 (.a(net_r[666]), .q(net_w[660]), .m(net_w[661]));
LSmitll_SPLITT_v2p1_optimized SC_474 (.a(net_r[667]), .q(net_w[662]), .m(net_w[663]));
LSmitll_SPLITT_v2p1_optimized SC_475 (.a(net_r[668]), .q(net_w[664]), .m(net_w[665]));
LSmitll_SPLITT_v2p1_optimized SC_476 (.a(net_r[669]), .q(net_w[666]), .m(net_w[667]));
LSmitll_SPLITT_v2p1_optimized SC_477 (.a(net_r[670]), .q(net_w[668]), .m());
LSmitll_SPLITT_v2p1_optimized SC_478 (.a(net_r[817]), .q(net_w[669]), .m(net_w[670]));
LSmitll_SPLITT_v2p1_optimized SC_479 (.a(net_r[682]), .q(net_w[671]), .m(net_w[672]));
LSmitll_SPLITT_v2p1_optimized SC_480 (.a(net_r[683]), .q(net_w[673]), .m(net_w[674]));
LSmitll_SPLITT_v2p1_optimized SC_481 (.a(net_r[684]), .q(net_w[675]), .m(net_w[676]));
LSmitll_SPLITT_v2p1_optimized SC_482 (.a(net_r[686]), .q(net_w[677]), .m(net_w[678]));
LSmitll_SPLITT_v2p1_optimized SC_483 (.a(net_r[687]), .q(net_w[679]), .m(net_w[680]));
LSmitll_SPLITT_v2p1_optimized SC_484 (.a(net_r[685]), .q(net_w[681]), .m());
LSmitll_SPLITT_v2p1_optimized SC_485 (.a(net_r[688]), .q(net_w[682]), .m(net_w[683]));
LSmitll_SPLITT_v2p1_optimized SC_486 (.a(net_r[689]), .q(net_w[684]), .m(net_w[685]));
LSmitll_SPLITT_v2p1_optimized SC_487 (.a(net_r[690]), .q(net_w[686]), .m(net_w[687]));
LSmitll_SPLITT_v2p1_optimized SC_488 (.a(net_r[691]), .q(net_w[688]), .m(net_w[689]));
LSmitll_SPLITT_v2p1_optimized SC_489 (.a(net_r[692]), .q(net_w[690]), .m());
LSmitll_SPLITT_v2p1_optimized SC_490 (.a(net_r[818]), .q(net_w[691]), .m(net_w[692]));
LSmitll_SPLITT_v2p1_optimized SC_491 (.a(net_r[703]), .q(net_w[693]), .m(net_w[694]));
LSmitll_SPLITT_v2p1_optimized SC_492 (.a(net_r[704]), .q(net_w[695]), .m(net_w[696]));
LSmitll_SPLITT_v2p1_optimized SC_493 (.a(net_r[705]), .q(net_w[697]), .m(net_w[698]));
LSmitll_SPLITT_v2p1_optimized SC_494 (.a(net_r[706]), .q(net_w[699]), .m(net_w[700]));
LSmitll_SPLITT_v2p1_optimized SC_495 (.a(net_r[707]), .q(net_w[701]), .m(net_w[702]));
LSmitll_SPLITT_v2p1_optimized SC_496 (.a(net_r[708]), .q(net_w[703]), .m(net_w[704]));
LSmitll_SPLITT_v2p1_optimized SC_497 (.a(net_r[710]), .q(net_w[705]), .m(net_w[706]));
LSmitll_SPLITT_v2p1_optimized SC_498 (.a(net_r[709]), .q(net_w[707]), .m());
LSmitll_SPLITT_v2p1_optimized SC_499 (.a(net_r[711]), .q(net_w[708]), .m(net_w[709]));
LSmitll_SPLITT_v2p1_optimized SC_500 (.a(net_r[712]), .q(net_w[710]), .m());
LSmitll_SPLITT_v2p1_optimized SC_501 (.a(net_r[819]), .q(net_w[711]), .m(net_w[712]));
LSmitll_SPLITT_v2p1_optimized SC_502 (.a(net_r[722]), .q(net_w[713]), .m(net_w[714]));
LSmitll_SPLITT_v2p1_optimized SC_503 (.a(net_r[723]), .q(net_w[715]), .m(net_w[716]));
LSmitll_SPLITT_v2p1_optimized SC_504 (.a(net_r[724]), .q(net_w[717]), .m(net_w[718]));
LSmitll_SPLITT_v2p1_optimized SC_505 (.a(net_r[726]), .q(net_w[719]), .m(net_w[720]));
LSmitll_SPLITT_v2p1_optimized SC_506 (.a(net_r[725]), .q(net_w[721]), .m());
LSmitll_SPLITT_v2p1_optimized SC_507 (.a(net_r[727]), .q(net_w[722]), .m(net_w[723]));
LSmitll_SPLITT_v2p1_optimized SC_508 (.a(net_r[729]), .q(net_w[724]), .m(net_w[725]));
LSmitll_SPLITT_v2p1_optimized SC_509 (.a(net_r[728]), .q(net_w[726]), .m());
LSmitll_SPLITT_v2p1_optimized SC_510 (.a(net_r[731]), .q(net_w[727]), .m(net_w[728]));
LSmitll_SPLITT_v2p1_optimized SC_511 (.a(net_r[730]), .q(net_w[729]), .m());
LSmitll_SPLITT_v2p1_optimized SC_512 (.a(net_r[820]), .q(net_w[730]), .m(net_w[731]));
LSmitll_SPLITT_v2p1_optimized SC_513 (.a(net_r[739]), .q(net_w[732]), .m(net_w[733]));
LSmitll_SPLITT_v2p1_optimized SC_514 (.a(net_r[740]), .q(net_w[734]), .m(net_w[735]));
LSmitll_SPLITT_v2p1_optimized SC_515 (.a(net_r[742]), .q(net_w[736]), .m(net_w[737]));
LSmitll_SPLITT_v2p1_optimized SC_516 (.a(net_r[741]), .q(net_w[738]), .m());
LSmitll_SPLITT_v2p1_optimized SC_517 (.a(net_r[743]), .q(net_w[739]), .m(net_w[740]));
LSmitll_SPLITT_v2p1_optimized SC_518 (.a(net_r[744]), .q(net_w[741]), .m(net_w[742]));
LSmitll_SPLITT_v2p1_optimized SC_519 (.a(net_r[745]), .q(net_w[743]), .m(net_w[744]));
LSmitll_SPLITT_v2p1_optimized SC_520 (.a(net_r[821]), .q(net_w[745]), .m());
LSmitll_SPLITT_v2p1_optimized SC_521 (.a(net_r[754]), .q(net_w[746]), .m(net_w[747]));
LSmitll_SPLITT_v2p1_optimized SC_522 (.a(net_r[755]), .q(net_w[748]), .m(net_w[749]));
LSmitll_SPLITT_v2p1_optimized SC_523 (.a(net_r[756]), .q(net_w[750]), .m(net_w[751]));
LSmitll_SPLITT_v2p1_optimized SC_524 (.a(net_r[757]), .q(net_w[752]), .m(net_w[753]));
LSmitll_SPLITT_v2p1_optimized SC_525 (.a(net_r[758]), .q(net_w[754]), .m(net_w[755]));
LSmitll_SPLITT_v2p1_optimized SC_526 (.a(net_r[759]), .q(net_w[756]), .m(net_w[757]));
LSmitll_SPLITT_v2p1_optimized SC_527 (.a(net_r[760]), .q(net_w[758]), .m(net_w[759]));
LSmitll_SPLITT_v2p1_optimized SC_528 (.a(net_r[822]), .q(net_w[760]), .m());
LSmitll_SPLITT_v2p1_optimized SC_529 (.a(net_r[768]), .q(net_w[761]), .m(net_w[762]));
LSmitll_SPLITT_v2p1_optimized SC_530 (.a(net_r[769]), .q(net_w[763]), .m(net_w[764]));
LSmitll_SPLITT_v2p1_optimized SC_531 (.a(net_r[771]), .q(net_w[765]), .m(net_w[766]));
LSmitll_SPLITT_v2p1_optimized SC_532 (.a(net_r[770]), .q(net_w[767]), .m());
LSmitll_SPLITT_v2p1_optimized SC_533 (.a(net_r[772]), .q(net_w[768]), .m(net_w[769]));
LSmitll_SPLITT_v2p1_optimized SC_534 (.a(net_r[773]), .q(net_w[770]), .m(net_w[771]));
LSmitll_SPLITT_v2p1_optimized SC_535 (.a(net_r[774]), .q(net_w[772]), .m(net_w[773]));
LSmitll_SPLITT_v2p1_optimized SC_536 (.a(net_r[823]), .q(net_w[774]), .m());
LSmitll_SPLITT_v2p1_optimized SC_537 (.a(net_r[780]), .q(net_w[775]), .m(net_w[776]));
LSmitll_SPLITT_v2p1_optimized SC_538 (.a(net_r[781]), .q(net_w[777]), .m(net_w[778]));
LSmitll_SPLITT_v2p1_optimized SC_539 (.a(net_r[782]), .q(net_w[779]), .m());
LSmitll_SPLITT_v2p1_optimized SC_540 (.a(net_r[783]), .q(net_w[780]), .m(net_w[781]));
LSmitll_SPLITT_v2p1_optimized SC_541 (.a(net_r[784]), .q(net_w[782]), .m());
LSmitll_SPLITT_v2p1_optimized SC_542 (.a(net_r[785]), .q(net_w[783]), .m(net_w[784]));
LSmitll_SPLITT_v2p1_optimized SC_543 (.a(net_r[824]), .q(net_w[785]), .m());
LSmitll_SPLITT_v2p1_optimized SC_544 (.a(net_r[789]), .q(net_w[786]), .m(net_w[787]));
LSmitll_SPLITT_v2p1_optimized SC_545 (.a(net_r[790]), .q(net_w[788]), .m());
LSmitll_SPLITT_v2p1_optimized SC_546 (.a(net_r[791]), .q(net_w[789]), .m(net_w[790]));
LSmitll_SPLITT_v2p1_optimized SC_547 (.a(net_r[792]), .q(net_w[791]), .m());
LSmitll_SPLITT_v2p1_optimized SC_548 (.a(net_r[825]), .q(net_w[792]), .m());
LSmitll_SPLITT_v2p1_optimized SC_549 (.a(net_r[796]), .q(net_w[793]), .m(net_w[794]));
LSmitll_SPLITT_v2p1_optimized SC_550 (.a(net_r[797]), .q(net_w[795]), .m());
LSmitll_SPLITT_v2p1_optimized SC_551 (.a(net_r[798]), .q(net_w[796]), .m(net_w[797]));
LSmitll_SPLITT_v2p1_optimized SC_552 (.a(net_r[799]), .q(net_w[798]), .m());
LSmitll_SPLITT_v2p1_optimized SC_553 (.a(net_r[826]), .q(net_w[799]), .m());
LSmitll_SPLITT_v2p1_optimized SC_554 (.a(net_r[332]), .q(net_w[800]), .m(net_w[801]));
LSmitll_SPLITT_v2p1_optimized SC_555 (.a(net_r[800]), .q(net_w[802]), .m(net_w[803]));
LSmitll_SPLITT_v2p1_optimized SC_556 (.a(net_r[801]), .q(net_w[804]), .m(net_w[805]));
LSmitll_SPLITT_v2p1_optimized SC_557 (.a(net_r[802]), .q(net_w[806]), .m(net_w[807]));
LSmitll_SPLITT_v2p1_optimized SC_558 (.a(net_r[803]), .q(net_w[808]), .m(net_w[809]));
LSmitll_SPLITT_v2p1_optimized SC_559 (.a(net_r[804]), .q(net_w[810]), .m(net_w[811]));
LSmitll_SPLITT_v2p1_optimized SC_560 (.a(net_r[805]), .q(net_w[812]), .m(net_w[813]));
LSmitll_SPLITT_v2p1_optimized SC_561 (.a(net_r[806]), .q(net_w[814]), .m(net_w[815]));
LSmitll_SPLITT_v2p1_optimized SC_562 (.a(net_r[807]), .q(net_w[816]), .m(net_w[817]));
LSmitll_SPLITT_v2p1_optimized SC_563 (.a(net_r[808]), .q(net_w[818]), .m(net_w[819]));
LSmitll_SPLITT_v2p1_optimized SC_564 (.a(net_r[809]), .q(net_w[820]), .m(net_w[821]));
LSmitll_SPLITT_v2p1_optimized SC_565 (.a(net_r[810]), .q(net_w[822]), .m(net_w[823]));
LSmitll_SPLITT_v2p1_optimized SC_566 (.a(net_r[811]), .q(net_w[824]), .m(net_w[825]));
LSmitll_SPLITT_v2p1_optimized SC_567 (.a(net_r[812]), .q(net_w[826]), .m());
LSmitll_SPLITT_v2p1_optimized SC_568 (.a(net_r[813]), .q(), .m());
endmodule