`include "data/modules/LSmitll_XORT_v2p1_selfcontained.v"
`include "data/modules/LSmitll_AND2T_v2p1_selfcontained.v"
`include "data/modules/LSmitll_SPLITT_v2p1_selfcontained.v"
`include "data/modules/LSmitll_OR2T_v2p1_selfcontained.v"
`include "data/modules/LSmitll_DFFT_v2p1_selfcontained.v"
`timescale 1ps/100fs
module KSA4 (
	A0,
	B0,
	SUM0,
	SUM1,
	SUM2,
	SUM3,
	COUT,
	A1,
	A2,
	A3,
	B1,
	B2,
	B3,
	CIN,
	clk
);
input
	A0,B0,A1,A2,A3,B1,B2,B3,CIN,clk;

output
	SUM0,SUM1,SUM2,SUM3,COUT;

reg  [252:0] net_r = 0;
wire [252:0] net_w;
assign net_w[1] = A0;
assign net_w[5] = B0;
assign net_w[31] = A1;
assign net_w[35] = A2;
assign net_w[41] = A3;
assign net_w[43] = B1;
assign net_w[47] = B2;
assign net_w[53] = B3;
assign net_w[54] = CIN;
assign net_w[107] = clk;
assign SUM0 = net_r[25];
assign SUM1 = net_r[26];
assign SUM2 = net_r[27];
assign SUM3 = net_r[28];
assign COUT = net_r[29];
always @(posedge net_w[1] or negedge net_w[1]) begin
	#1.40097 net_r[1] <= net_w[1];
end
always @(posedge net_w[2] or negedge net_w[2]) begin
	#0.500346 net_r[2] <= net_w[2];
end
always @(posedge net_w[3] or negedge net_w[3]) begin
	#0.700485 net_r[3] <= net_w[3];
end
always @(posedge net_w[4] or negedge net_w[4]) begin
	#0.800554 net_r[4] <= net_w[4];
end
always @(posedge net_w[5] or negedge net_w[5]) begin
	#1.10076 net_r[5] <= net_w[5];
end
always @(posedge net_w[6] or negedge net_w[6]) begin
	#0.500346 net_r[6] <= net_w[6];
end
always @(posedge net_w[7] or negedge net_w[7]) begin
	#0.800554 net_r[7] <= net_w[7];
end
always @(posedge net_w[8] or negedge net_w[8]) begin
	#0.500346 net_r[8] <= net_w[8];
end
always @(posedge net_w[9] or negedge net_w[9]) begin
	#1.40097 net_r[9] <= net_w[9];
end
always @(posedge net_w[10] or negedge net_w[10]) begin
	#0.500346 net_r[10] <= net_w[10];
end
always @(posedge net_w[11] or negedge net_w[11]) begin
	#2.70187 net_r[11] <= net_w[11];
end
always @(posedge net_w[12] or negedge net_w[12]) begin
	#0.500346 net_r[12] <= net_w[12];
end
always @(posedge net_w[13] or negedge net_w[13]) begin
	#2.00138 net_r[13] <= net_w[13];
end
always @(posedge net_w[14] or negedge net_w[14]) begin
	#0.500346 net_r[14] <= net_w[14];
end
always @(posedge net_w[15] or negedge net_w[15]) begin
	#5.10353 net_r[15] <= net_w[15];
end
always @(posedge net_w[16] or negedge net_w[16]) begin
	#2.00138 net_r[16] <= net_w[16];
end
always @(posedge net_w[17] or negedge net_w[17]) begin
	#0.800554 net_r[17] <= net_w[17];
end
always @(posedge net_w[18] or negedge net_w[18]) begin
	#1.60111 net_r[18] <= net_w[18];
end
always @(posedge net_w[19] or negedge net_w[19]) begin
	#5.2036 net_r[19] <= net_w[19];
end
always @(posedge net_w[20] or negedge net_w[20]) begin
	#0.900623 net_r[20] <= net_w[20];
end
always @(posedge net_w[21] or negedge net_w[21]) begin
	#2.20152 net_r[21] <= net_w[21];
end
always @(posedge net_w[22] or negedge net_w[22]) begin
	#0.500346 net_r[22] <= net_w[22];
end
always @(posedge net_w[23] or negedge net_w[23]) begin
	#8.60595 net_r[23] <= net_w[23];
end
always @(posedge net_w[24] or negedge net_w[24]) begin
	#2.90201 net_r[24] <= net_w[24];
end
always @(posedge net_w[25] or negedge net_w[25]) begin
	#5.80402 net_r[25] <= net_w[25];
end
always @(posedge net_w[26] or negedge net_w[26]) begin
	#3.50242 net_r[26] <= net_w[26];
end
always @(posedge net_w[27] or negedge net_w[27]) begin
	#3.20222 net_r[27] <= net_w[27];
end
always @(posedge net_w[28] or negedge net_w[28]) begin
	#3.10215 net_r[28] <= net_w[28];
end
always @(posedge net_w[29] or negedge net_w[29]) begin
	#1.50104 net_r[29] <= net_w[29];
end
always @(posedge net_w[30] or negedge net_w[30]) begin
	#2.00138 net_r[30] <= net_w[30];
end
always @(posedge net_w[31] or negedge net_w[31]) begin
	#1.90132 net_r[31] <= net_w[31];
end
always @(posedge net_w[32] or negedge net_w[32]) begin
	#2.20152 net_r[32] <= net_w[32];
end
always @(posedge net_w[33] or negedge net_w[33]) begin
	#1.10076 net_r[33] <= net_w[33];
end
always @(posedge net_w[34] or negedge net_w[34]) begin
	#2.00138 net_r[34] <= net_w[34];
end
always @(posedge net_w[35] or negedge net_w[35]) begin
	#1.80125 net_r[35] <= net_w[35];
end
always @(posedge net_w[36] or negedge net_w[36]) begin
	#2.00138 net_r[36] <= net_w[36];
end
always @(posedge net_w[37] or negedge net_w[37]) begin
	#1.20083 net_r[37] <= net_w[37];
end
always @(posedge net_w[38] or negedge net_w[38]) begin
	#2.00138 net_r[38] <= net_w[38];
end
always @(posedge net_w[39] or negedge net_w[39]) begin
	#1.00069 net_r[39] <= net_w[39];
end
always @(posedge net_w[40] or negedge net_w[40]) begin
	#2.10145 net_r[40] <= net_w[40];
end
always @(posedge net_w[41] or negedge net_w[41]) begin
	#1.70118 net_r[41] <= net_w[41];
end
always @(posedge net_w[42] or negedge net_w[42]) begin
	#1.70118 net_r[42] <= net_w[42];
end
always @(posedge net_w[43] or negedge net_w[43]) begin
	#1.70118 net_r[43] <= net_w[43];
end
always @(posedge net_w[44] or negedge net_w[44]) begin
	#1.90132 net_r[44] <= net_w[44];
end
always @(posedge net_w[45] or negedge net_w[45]) begin
	#1.00069 net_r[45] <= net_w[45];
end
always @(posedge net_w[46] or negedge net_w[46]) begin
	#1.70118 net_r[46] <= net_w[46];
end
always @(posedge net_w[47] or negedge net_w[47]) begin
	#1.60111 net_r[47] <= net_w[47];
end
always @(posedge net_w[48] or negedge net_w[48]) begin
	#2.30159 net_r[48] <= net_w[48];
end
always @(posedge net_w[49] or negedge net_w[49]) begin
	#1.40097 net_r[49] <= net_w[49];
end
always @(posedge net_w[50] or negedge net_w[50]) begin
	#2.00138 net_r[50] <= net_w[50];
end
always @(posedge net_w[51] or negedge net_w[51]) begin
	#0.900623 net_r[51] <= net_w[51];
end
always @(posedge net_w[52] or negedge net_w[52]) begin
	#1.80125 net_r[52] <= net_w[52];
end
always @(posedge net_w[53] or negedge net_w[53]) begin
	#1.40097 net_r[53] <= net_w[53];
end
always @(posedge net_w[54] or negedge net_w[54]) begin
	#1.3009 net_r[54] <= net_w[54];
end
always @(posedge net_w[55] or negedge net_w[55]) begin
	#1.10076 net_r[55] <= net_w[55];
end
always @(posedge net_w[56] or negedge net_w[56]) begin
	#1.20083 net_r[56] <= net_w[56];
end
always @(posedge net_w[57] or negedge net_w[57]) begin
	#1.40097 net_r[57] <= net_w[57];
end
always @(posedge net_w[58] or negedge net_w[58]) begin
	#1.40097 net_r[58] <= net_w[58];
end
always @(posedge net_w[59] or negedge net_w[59]) begin
	#1.3009 net_r[59] <= net_w[59];
end
always @(posedge net_w[60] or negedge net_w[60]) begin
	#2.90201 net_r[60] <= net_w[60];
end
always @(posedge net_w[61] or negedge net_w[61]) begin
	#1.40097 net_r[61] <= net_w[61];
end
always @(posedge net_w[62] or negedge net_w[62]) begin
	#2.6018 net_r[62] <= net_w[62];
end
always @(posedge net_w[63] or negedge net_w[63]) begin
	#0.900623 net_r[63] <= net_w[63];
end
always @(posedge net_w[64] or negedge net_w[64]) begin
	#2.50173 net_r[64] <= net_w[64];
end
always @(posedge net_w[65] or negedge net_w[65]) begin
	#1.00069 net_r[65] <= net_w[65];
end
always @(posedge net_w[66] or negedge net_w[66]) begin
	#3.9027 net_r[66] <= net_w[66];
end
always @(posedge net_w[67] or negedge net_w[67]) begin
	#1.10076 net_r[67] <= net_w[67];
end
always @(posedge net_w[68] or negedge net_w[68]) begin
	#2.6018 net_r[68] <= net_w[68];
end
always @(posedge net_w[69] or negedge net_w[69]) begin
	#1.40097 net_r[69] <= net_w[69];
end
always @(posedge net_w[70] or negedge net_w[70]) begin
	#2.50173 net_r[70] <= net_w[70];
end
always @(posedge net_w[71] or negedge net_w[71]) begin
	#2.70187 net_r[71] <= net_w[71];
end
always @(posedge net_w[72] or negedge net_w[72]) begin
	#3.10215 net_r[72] <= net_w[72];
end
always @(posedge net_w[73] or negedge net_w[73]) begin
	#0.900623 net_r[73] <= net_w[73];
end
always @(posedge net_w[74] or negedge net_w[74]) begin
	#4.20291 net_r[74] <= net_w[74];
end
always @(posedge net_w[75] or negedge net_w[75]) begin
	#1.70118 net_r[75] <= net_w[75];
end
always @(posedge net_w[76] or negedge net_w[76]) begin
	#1.90132 net_r[76] <= net_w[76];
end
always @(posedge net_w[77] or negedge net_w[77]) begin
	#1.60111 net_r[77] <= net_w[77];
end
always @(posedge net_w[78] or negedge net_w[78]) begin
	#2.10145 net_r[78] <= net_w[78];
end
always @(posedge net_w[79] or negedge net_w[79]) begin
	#3.10215 net_r[79] <= net_w[79];
end
always @(posedge net_w[80] or negedge net_w[80]) begin
	#2.40166 net_r[80] <= net_w[80];
end
always @(posedge net_w[81] or negedge net_w[81]) begin
	#2.70187 net_r[81] <= net_w[81];
end
always @(posedge net_w[82] or negedge net_w[82]) begin
	#1.80125 net_r[82] <= net_w[82];
end
always @(posedge net_w[83] or negedge net_w[83]) begin
	#5.40374 net_r[83] <= net_w[83];
end
always @(posedge net_w[84] or negedge net_w[84]) begin
	#3.30228 net_r[84] <= net_w[84];
end
always @(posedge net_w[85] or negedge net_w[85]) begin
	#4.70325 net_r[85] <= net_w[85];
end
always @(posedge net_w[86] or negedge net_w[86]) begin
	#2.70187 net_r[86] <= net_w[86];
end
always @(posedge net_w[87] or negedge net_w[87]) begin
	#5.30367 net_r[87] <= net_w[87];
end
always @(posedge net_w[88] or negedge net_w[88]) begin
	#2.90201 net_r[88] <= net_w[88];
end
always @(posedge net_w[89] or negedge net_w[89]) begin
	#4.00277 net_r[89] <= net_w[89];
end
always @(posedge net_w[90] or negedge net_w[90]) begin
	#1.40097 net_r[90] <= net_w[90];
end
always @(posedge net_w[91] or negedge net_w[91]) begin
	#9.1063 net_r[91] <= net_w[91];
end
always @(posedge net_w[92] or negedge net_w[92]) begin
	#8.70602 net_r[92] <= net_w[92];
end
always @(posedge net_w[93] or negedge net_w[93]) begin
	#2.40166 net_r[93] <= net_w[93];
end
always @(posedge net_w[94] or negedge net_w[94]) begin
	#1.90132 net_r[94] <= net_w[94];
end
always @(posedge net_w[95] or negedge net_w[95]) begin
	#0.800554 net_r[95] <= net_w[95];
end
always @(posedge net_w[96] or negedge net_w[96]) begin
	#2.20152 net_r[96] <= net_w[96];
end
always @(posedge net_w[97] or negedge net_w[97]) begin
	#3.30228 net_r[97] <= net_w[97];
end
always @(posedge net_w[98] or negedge net_w[98]) begin
	#3.20222 net_r[98] <= net_w[98];
end
always @(posedge net_w[99] or negedge net_w[99]) begin
	#1.40097 net_r[99] <= net_w[99];
end
always @(posedge net_w[100] or negedge net_w[100]) begin
	#3.00208 net_r[100] <= net_w[100];
end
always @(posedge net_w[101] or negedge net_w[101]) begin
	#4.40305 net_r[101] <= net_w[101];
end
always @(posedge net_w[102] or negedge net_w[102]) begin
	#5.70395 net_r[102] <= net_w[102];
end
always @(posedge net_w[103] or negedge net_w[103]) begin
	#2.20152 net_r[103] <= net_w[103];
end
always @(posedge net_w[104] or negedge net_w[104]) begin
	#1.00069 net_r[104] <= net_w[104];
end
always @(posedge net_w[105] or negedge net_w[105]) begin
	#6.10422 net_r[105] <= net_w[105];
end
always @(posedge net_w[106] or negedge net_w[106]) begin
	#5.40374 net_r[106] <= net_w[106];
end
always @(posedge net_w[107] or negedge net_w[107]) begin
	#8.60595 net_r[107] <= net_w[107];
end
always @(posedge net_w[108] or negedge net_w[108]) begin
	#1.50104 net_r[108] <= net_w[108];
end
always @(posedge net_w[109] or negedge net_w[109]) begin
	#2.10145 net_r[109] <= net_w[109];
end
always @(posedge net_w[110] or negedge net_w[110]) begin
	#0.400277 net_r[110] <= net_w[110];
end
always @(posedge net_w[111] or negedge net_w[111]) begin
	#1.90132 net_r[111] <= net_w[111];
end
always @(posedge net_w[112] or negedge net_w[112]) begin
	#0.400277 net_r[112] <= net_w[112];
end
always @(posedge net_w[113] or negedge net_w[113]) begin
	#1.70118 net_r[113] <= net_w[113];
end
always @(posedge net_w[114] or negedge net_w[114]) begin
	#0.600415 net_r[114] <= net_w[114];
end
always @(posedge net_w[115] or negedge net_w[115]) begin
	#0.900623 net_r[115] <= net_w[115];
end
always @(posedge net_w[116] or negedge net_w[116]) begin
	#1.50104 net_r[116] <= net_w[116];
end
always @(posedge net_w[117] or negedge net_w[117]) begin
	#0.700485 net_r[117] <= net_w[117];
end
always @(posedge net_w[118] or negedge net_w[118]) begin
	#1.50104 net_r[118] <= net_w[118];
end
always @(posedge net_w[119] or negedge net_w[119]) begin
	#0.500346 net_r[119] <= net_w[119];
end
always @(posedge net_w[120] or negedge net_w[120]) begin
	#1.40097 net_r[120] <= net_w[120];
end
always @(posedge net_w[121] or negedge net_w[121]) begin
	#0.500346 net_r[121] <= net_w[121];
end
always @(posedge net_w[122] or negedge net_w[122]) begin
	#1.60111 net_r[122] <= net_w[122];
end
always @(posedge net_w[123] or negedge net_w[123]) begin
	#1.50104 net_r[123] <= net_w[123];
end
always @(posedge net_w[124] or negedge net_w[124]) begin
	#2.40166 net_r[124] <= net_w[124];
end
always @(posedge net_w[125] or negedge net_w[125]) begin
	#0.400277 net_r[125] <= net_w[125];
end
always @(posedge net_w[126] or negedge net_w[126]) begin
	#2.10145 net_r[126] <= net_w[126];
end
always @(posedge net_w[127] or negedge net_w[127]) begin
	#2.10145 net_r[127] <= net_w[127];
end
always @(posedge net_w[128] or negedge net_w[128]) begin
	#1.20083 net_r[128] <= net_w[128];
end
always @(posedge net_w[129] or negedge net_w[129]) begin
	#1.50104 net_r[129] <= net_w[129];
end
always @(posedge net_w[130] or negedge net_w[130]) begin
	#0.600415 net_r[130] <= net_w[130];
end
always @(posedge net_w[131] or negedge net_w[131]) begin
	#1.3009 net_r[131] <= net_w[131];
end
always @(posedge net_w[132] or negedge net_w[132]) begin
	#1.60111 net_r[132] <= net_w[132];
end
always @(posedge net_w[133] or negedge net_w[133]) begin
	#1.00069 net_r[133] <= net_w[133];
end
always @(posedge net_w[134] or negedge net_w[134]) begin
	#1.3009 net_r[134] <= net_w[134];
end
always @(posedge net_w[135] or negedge net_w[135]) begin
	#0.700485 net_r[135] <= net_w[135];
end
always @(posedge net_w[136] or negedge net_w[136]) begin
	#1.80125 net_r[136] <= net_w[136];
end
always @(posedge net_w[137] or negedge net_w[137]) begin
	#0.400277 net_r[137] <= net_w[137];
end
always @(posedge net_w[138] or negedge net_w[138]) begin
	#2.10145 net_r[138] <= net_w[138];
end
always @(posedge net_w[139] or negedge net_w[139]) begin
	#1.90132 net_r[139] <= net_w[139];
end
always @(posedge net_w[140] or negedge net_w[140]) begin
	#2.50173 net_r[140] <= net_w[140];
end
always @(posedge net_w[141] or negedge net_w[141]) begin
	#1.00069 net_r[141] <= net_w[141];
end
always @(posedge net_w[142] or negedge net_w[142]) begin
	#1.40097 net_r[142] <= net_w[142];
end
always @(posedge net_w[143] or negedge net_w[143]) begin
	#2.50173 net_r[143] <= net_w[143];
end
always @(posedge net_w[144] or negedge net_w[144]) begin
	#0.900623 net_r[144] <= net_w[144];
end
always @(posedge net_w[145] or negedge net_w[145]) begin
	#1.70118 net_r[145] <= net_w[145];
end
always @(posedge net_w[146] or negedge net_w[146]) begin
	#2.00138 net_r[146] <= net_w[146];
end
always @(posedge net_w[147] or negedge net_w[147]) begin
	#0.500346 net_r[147] <= net_w[147];
end
always @(posedge net_w[148] or negedge net_w[148]) begin
	#2.40166 net_r[148] <= net_w[148];
end
always @(posedge net_w[149] or negedge net_w[149]) begin
	#0.500346 net_r[149] <= net_w[149];
end
always @(posedge net_w[150] or negedge net_w[150]) begin
	#2.20152 net_r[150] <= net_w[150];
end
always @(posedge net_w[151] or negedge net_w[151]) begin
	#1.00069 net_r[151] <= net_w[151];
end
always @(posedge net_w[152] or negedge net_w[152]) begin
	#1.3009 net_r[152] <= net_w[152];
end
always @(posedge net_w[153] or negedge net_w[153]) begin
	#2.50173 net_r[153] <= net_w[153];
end
always @(posedge net_w[154] or negedge net_w[154]) begin
	#1.20083 net_r[154] <= net_w[154];
end
always @(posedge net_w[155] or negedge net_w[155]) begin
	#2.40166 net_r[155] <= net_w[155];
end
always @(posedge net_w[156] or negedge net_w[156]) begin
	#0.600415 net_r[156] <= net_w[156];
end
always @(posedge net_w[157] or negedge net_w[157]) begin
	#1.40097 net_r[157] <= net_w[157];
end
always @(posedge net_w[158] or negedge net_w[158]) begin
	#1.3009 net_r[158] <= net_w[158];
end
always @(posedge net_w[159] or negedge net_w[159]) begin
	#0.800554 net_r[159] <= net_w[159];
end
always @(posedge net_w[160] or negedge net_w[160]) begin
	#1.10076 net_r[160] <= net_w[160];
end
always @(posedge net_w[161] or negedge net_w[161]) begin
	#1.70118 net_r[161] <= net_w[161];
end
always @(posedge net_w[162] or negedge net_w[162]) begin
	#2.40166 net_r[162] <= net_w[162];
end
always @(posedge net_w[163] or negedge net_w[163]) begin
	#1.00069 net_r[163] <= net_w[163];
end
always @(posedge net_w[164] or negedge net_w[164]) begin
	#1.60111 net_r[164] <= net_w[164];
end
always @(posedge net_w[165] or negedge net_w[165]) begin
	#0.600415 net_r[165] <= net_w[165];
end
always @(posedge net_w[166] or negedge net_w[166]) begin
	#3.20222 net_r[166] <= net_w[166];
end
always @(posedge net_w[167] or negedge net_w[167]) begin
	#1.3009 net_r[167] <= net_w[167];
end
always @(posedge net_w[168] or negedge net_w[168]) begin
	#2.80194 net_r[168] <= net_w[168];
end
always @(posedge net_w[169] or negedge net_w[169]) begin
	#1.60111 net_r[169] <= net_w[169];
end
always @(posedge net_w[170] or negedge net_w[170]) begin
	#2.20152 net_r[170] <= net_w[170];
end
always @(posedge net_w[171] or negedge net_w[171]) begin
	#2.20152 net_r[171] <= net_w[171];
end
always @(posedge net_w[172] or negedge net_w[172]) begin
	#2.30159 net_r[172] <= net_w[172];
end
always @(posedge net_w[173] or negedge net_w[173]) begin
	#1.10076 net_r[173] <= net_w[173];
end
always @(posedge net_w[174] or negedge net_w[174]) begin
	#0.700485 net_r[174] <= net_w[174];
end
always @(posedge net_w[175] or negedge net_w[175]) begin
	#0.900623 net_r[175] <= net_w[175];
end
always @(posedge net_w[176] or negedge net_w[176]) begin
	#0.700485 net_r[176] <= net_w[176];
end
always @(posedge net_w[177] or negedge net_w[177]) begin
	#0.900623 net_r[177] <= net_w[177];
end
always @(posedge net_w[178] or negedge net_w[178]) begin
	#0.700485 net_r[178] <= net_w[178];
end
always @(posedge net_w[179] or negedge net_w[179]) begin
	#0.900623 net_r[179] <= net_w[179];
end
always @(posedge net_w[180] or negedge net_w[180]) begin
	#0.700485 net_r[180] <= net_w[180];
end
always @(posedge net_w[181] or negedge net_w[181]) begin
	#1.60111 net_r[181] <= net_w[181];
end
always @(posedge net_w[182] or negedge net_w[182]) begin
	#1.40097 net_r[182] <= net_w[182];
end
always @(posedge net_w[183] or negedge net_w[183]) begin
	#1.80125 net_r[183] <= net_w[183];
end
always @(posedge net_w[184] or negedge net_w[184]) begin
	#1.20083 net_r[184] <= net_w[184];
end
always @(posedge net_w[185] or negedge net_w[185]) begin
	#2.80194 net_r[185] <= net_w[185];
end
always @(posedge net_w[186] or negedge net_w[186]) begin
	#2.40166 net_r[186] <= net_w[186];
end
always @(posedge net_w[187] or negedge net_w[187]) begin
	#2.10145 net_r[187] <= net_w[187];
end
always @(posedge net_w[188] or negedge net_w[188]) begin
	#0.700485 net_r[188] <= net_w[188];
end
always @(posedge net_w[189] or negedge net_w[189]) begin
	#0.900623 net_r[189] <= net_w[189];
end
always @(posedge net_w[190] or negedge net_w[190]) begin
	#1.3009 net_r[190] <= net_w[190];
end
always @(posedge net_w[191] or negedge net_w[191]) begin
	#0.900623 net_r[191] <= net_w[191];
end
always @(posedge net_w[192] or negedge net_w[192]) begin
	#1.3009 net_r[192] <= net_w[192];
end
always @(posedge net_w[193] or negedge net_w[193]) begin
	#3.50242 net_r[193] <= net_w[193];
end
always @(posedge net_w[194] or negedge net_w[194]) begin
	#1.50104 net_r[194] <= net_w[194];
end
always @(posedge net_w[195] or negedge net_w[195]) begin
	#2.40166 net_r[195] <= net_w[195];
end
always @(posedge net_w[196] or negedge net_w[196]) begin
	#1.40097 net_r[196] <= net_w[196];
end
always @(posedge net_w[197] or negedge net_w[197]) begin
	#0.700485 net_r[197] <= net_w[197];
end
always @(posedge net_w[198] or negedge net_w[198]) begin
	#3.20222 net_r[198] <= net_w[198];
end
always @(posedge net_w[199] or negedge net_w[199]) begin
	#2.00138 net_r[199] <= net_w[199];
end
always @(posedge net_w[200] or negedge net_w[200]) begin
	#1.50104 net_r[200] <= net_w[200];
end
always @(posedge net_w[201] or negedge net_w[201]) begin
	#0.800554 net_r[201] <= net_w[201];
end
always @(posedge net_w[202] or negedge net_w[202]) begin
	#1.10076 net_r[202] <= net_w[202];
end
always @(posedge net_w[203] or negedge net_w[203]) begin
	#1.50104 net_r[203] <= net_w[203];
end
always @(posedge net_w[204] or negedge net_w[204]) begin
	#1.80125 net_r[204] <= net_w[204];
end
always @(posedge net_w[205] or negedge net_w[205]) begin
	#1.70118 net_r[205] <= net_w[205];
end
always @(posedge net_w[206] or negedge net_w[206]) begin
	#3.10215 net_r[206] <= net_w[206];
end
always @(posedge net_w[207] or negedge net_w[207]) begin
	#2.6018 net_r[207] <= net_w[207];
end
always @(posedge net_w[208] or negedge net_w[208]) begin
	#1.10076 net_r[208] <= net_w[208];
end
always @(posedge net_w[209] or negedge net_w[209]) begin
	#0.800554 net_r[209] <= net_w[209];
end
always @(posedge net_w[210] or negedge net_w[210]) begin
	#1.10076 net_r[210] <= net_w[210];
end
always @(posedge net_w[211] or negedge net_w[211]) begin
	#0.800554 net_r[211] <= net_w[211];
end
always @(posedge net_w[212] or negedge net_w[212]) begin
	#1.10076 net_r[212] <= net_w[212];
end
always @(posedge net_w[213] or negedge net_w[213]) begin
	#1.50104 net_r[213] <= net_w[213];
end
always @(posedge net_w[214] or negedge net_w[214]) begin
	#1.80125 net_r[214] <= net_w[214];
end
always @(posedge net_w[215] or negedge net_w[215]) begin
	#1.70118 net_r[215] <= net_w[215];
end
always @(posedge net_w[216] or negedge net_w[216]) begin
	#4.10284 net_r[216] <= net_w[216];
end
always @(posedge net_w[217] or negedge net_w[217]) begin
	#2.6018 net_r[217] <= net_w[217];
end
always @(posedge net_w[218] or negedge net_w[218]) begin
	#1.10076 net_r[218] <= net_w[218];
end
always @(posedge net_w[219] or negedge net_w[219]) begin
	#0.800554 net_r[219] <= net_w[219];
end
always @(posedge net_w[220] or negedge net_w[220]) begin
	#1.70118 net_r[220] <= net_w[220];
end
always @(posedge net_w[221] or negedge net_w[221]) begin
	#2.00138 net_r[221] <= net_w[221];
end
always @(posedge net_w[222] or negedge net_w[222]) begin
	#1.3009 net_r[222] <= net_w[222];
end
always @(posedge net_w[223] or negedge net_w[223]) begin
	#1.10076 net_r[223] <= net_w[223];
end
always @(posedge net_w[224] or negedge net_w[224]) begin
	#3.10215 net_r[224] <= net_w[224];
end
always @(posedge net_w[225] or negedge net_w[225]) begin
	#2.00138 net_r[225] <= net_w[225];
end
always @(posedge net_w[226] or negedge net_w[226]) begin
	#2.20152 net_r[226] <= net_w[226];
end
always @(posedge net_w[227] or negedge net_w[227]) begin
	#1.40097 net_r[227] <= net_w[227];
end
always @(posedge net_w[228] or negedge net_w[228]) begin
	#2.20152 net_r[228] <= net_w[228];
end
always @(posedge net_w[229] or negedge net_w[229]) begin
	#1.40097 net_r[229] <= net_w[229];
end
always @(posedge net_w[230] or negedge net_w[230]) begin
	#3.40235 net_r[230] <= net_w[230];
end
always @(posedge net_w[231] or negedge net_w[231]) begin
	#1.20083 net_r[231] <= net_w[231];
end
always @(posedge net_w[232] or negedge net_w[232]) begin
	#2.40166 net_r[232] <= net_w[232];
end
always @(posedge net_w[233] or negedge net_w[233]) begin
	#1.40097 net_r[233] <= net_w[233];
end
always @(posedge net_w[234] or negedge net_w[234]) begin
	#2.20152 net_r[234] <= net_w[234];
end
always @(posedge net_w[235] or negedge net_w[235]) begin
	#1.40097 net_r[235] <= net_w[235];
end
always @(posedge net_w[236] or negedge net_w[236]) begin
	#3.60249 net_r[236] <= net_w[236];
end
always @(posedge net_w[237] or negedge net_w[237]) begin
	#1.20083 net_r[237] <= net_w[237];
end
always @(posedge net_w[238] or negedge net_w[238]) begin
	#2.40166 net_r[238] <= net_w[238];
end
always @(posedge net_w[239] or negedge net_w[239]) begin
	#5.70395 net_r[239] <= net_w[239];
end
always @(posedge net_w[240] or negedge net_w[240]) begin
	#4.80332 net_r[240] <= net_w[240];
end
always @(posedge net_w[241] or negedge net_w[241]) begin
	#3.30228 net_r[241] <= net_w[241];
end
always @(posedge net_w[242] or negedge net_w[242]) begin
	#2.20152 net_r[242] <= net_w[242];
end
always @(posedge net_w[243] or negedge net_w[243]) begin
	#3.10215 net_r[243] <= net_w[243];
end
always @(posedge net_w[244] or negedge net_w[244]) begin
	#2.00138 net_r[244] <= net_w[244];
end
always @(posedge net_w[245] or negedge net_w[245]) begin
	#4.70325 net_r[245] <= net_w[245];
end
always @(posedge net_w[246] or negedge net_w[246]) begin
	#7.00485 net_r[246] <= net_w[246];
end
always @(posedge net_w[247] or negedge net_w[247]) begin
	#3.9027 net_r[247] <= net_w[247];
end
always @(posedge net_w[248] or negedge net_w[248]) begin
	#5.30367 net_r[248] <= net_w[248];
end
always @(posedge net_w[249] or negedge net_w[249]) begin
	#2.00138 net_r[249] <= net_w[249];
end
always @(posedge net_w[250] or negedge net_w[250]) begin
	#4.60318 net_r[250] <= net_w[250];
end
always @(posedge net_w[251] or negedge net_w[251]) begin
	#2.10145 net_r[251] <= net_w[251];
end
LSmitll_XORT_v2p1_optimized XOR2T_0 (.a(net_r[75]), .b(net_r[83]), .clk(net_r[108]), .q(net_w[10]));
LSmitll_XORT_v2p1_optimized XOR2T_1 (.a(net_r[91]), .b(net_r[93]), .clk(net_r[123]), .q(net_w[65]));
LSmitll_AND2T AND2T_2 (.a(net_r[76]), .b(net_r[84]), .clk(net_r[110]), .q(net_w[55]));
LSmitll_AND2T AND2T_3 (.a(net_r[92]), .b(net_r[94]), .clk(net_r[125]), .q(net_w[12]));
LSmitll_OR2T_v2p1_optimized OR2T_4 (.a(net_r[11]), .b(net_r[12]), .clk(net_r[138]), .q(net_w[13]));
LSmitll_XORT_v2p1_optimized XOR2T_5 (.a(net_r[77]), .b(net_r[85]), .clk(net_r[126]), .q(net_w[14]));
LSmitll_XORT_v2p1_optimized XOR2T_6 (.a(net_r[95]), .b(net_r[97]), .clk(net_r[148]), .q(net_w[70]));
LSmitll_AND2T AND2T_7 (.a(net_r[78]), .b(net_r[86]), .clk(net_r[128]), .q(net_w[56]));
LSmitll_AND2T AND2T_8 (.a(net_r[96]), .b(net_r[98]), .clk(net_r[150]), .q(net_w[16]));
LSmitll_OR2T_v2p1_optimized OR2T_9 (.a(net_r[15]), .b(net_r[16]), .clk(net_r[151]), .q(net_w[17]));
LSmitll_XORT_v2p1_optimized XOR2T_10 (.a(net_r[79]), .b(net_r[87]), .clk(net_r[139]), .q(net_w[18]));
LSmitll_XORT_v2p1_optimized XOR2T_11 (.a(net_r[99]), .b(net_r[101]), .clk(net_r[159]), .q(net_w[73]));
LSmitll_AND2T AND2T_12 (.a(net_r[80]), .b(net_r[88]), .clk(net_r[141]), .q(net_w[57]));
LSmitll_AND2T AND2T_13 (.a(net_r[100]), .b(net_r[102]), .clk(net_r[160]), .q(net_w[20]));
LSmitll_OR2T_v2p1_optimized OR2T_14 (.a(net_r[19]), .b(net_r[20]), .clk(net_r[167]), .q(net_w[21]));
LSmitll_XORT_v2p1_optimized XOR2T_15 (.a(net_r[81]), .b(net_r[89]), .clk(net_r[152]), .q(net_w[22]));
LSmitll_XORT_v2p1_optimized XOR2T_16 (.a(net_r[103]), .b(net_r[105]), .clk(net_r[170]), .q(net_w[74]));
LSmitll_AND2T AND2T_17 (.a(net_r[82]), .b(net_r[90]), .clk(net_r[154]), .q(net_w[58]));
LSmitll_AND2T AND2T_18 (.a(net_r[104]), .b(net_r[106]), .clk(net_r[172]), .q(net_w[24]));
LSmitll_OR2T_v2p1_optimized OR2T_19 (.a(net_r[23]), .b(net_r[24]), .clk(net_r[171]), .q(net_w[29]));
LSmitll_DFFT_v2p1_optimized DFF_34 (.a(net_r[30]), .clk(net_r[112]), .q(net_w[2]));
LSmitll_DFFT_v2p1_optimized DFF_35 (.a(net_r[31]), .clk(net_r[109]), .q(net_w[30]));
LSmitll_DFFT_v2p1_optimized DFF_36 (.a(net_r[32]), .clk(net_r[130]), .q(net_w[3]));
LSmitll_DFFT_v2p1_optimized DFF_37 (.a(net_r[33]), .clk(net_r[127]), .q(net_w[32]));
LSmitll_DFFT_v2p1_optimized DFF_38 (.a(net_r[34]), .clk(net_r[114]), .q(net_w[33]));
LSmitll_DFFT_v2p1_optimized DFF_39 (.a(net_r[35]), .clk(net_r[111]), .q(net_w[34]));
LSmitll_DFFT_v2p1_optimized DFF_40 (.a(net_r[36]), .clk(net_r[142]), .q(net_w[4]));
LSmitll_DFFT_v2p1_optimized DFF_41 (.a(net_r[37]), .clk(net_r[143]), .q(net_w[36]));
LSmitll_DFFT_v2p1_optimized DFF_42 (.a(net_r[38]), .clk(net_r[131]), .q(net_w[37]));
LSmitll_DFFT_v2p1_optimized DFF_43 (.a(net_r[39]), .clk(net_r[129]), .q(net_w[38]));
LSmitll_DFFT_v2p1_optimized DFF_44 (.a(net_r[40]), .clk(net_r[115]), .q(net_w[39]));
LSmitll_DFFT_v2p1_optimized DFF_45 (.a(net_r[41]), .clk(net_r[113]), .q(net_w[40]));
LSmitll_DFFT_v2p1_optimized DFF_46 (.a(net_r[42]), .clk(net_r[117]), .q(net_w[6]));
LSmitll_DFFT_v2p1_optimized DFF_47 (.a(net_r[43]), .clk(net_r[116]), .q(net_w[42]));
LSmitll_DFFT_v2p1_optimized DFF_48 (.a(net_r[44]), .clk(net_r[133]), .q(net_w[7]));
LSmitll_DFFT_v2p1_optimized DFF_49 (.a(net_r[45]), .clk(net_r[132]), .q(net_w[44]));
LSmitll_DFFT_v2p1_optimized DFF_50 (.a(net_r[46]), .clk(net_r[119]), .q(net_w[45]));
LSmitll_DFFT_v2p1_optimized DFF_51 (.a(net_r[47]), .clk(net_r[118]), .q(net_w[46]));
LSmitll_DFFT_v2p1_optimized DFF_52 (.a(net_r[48]), .clk(net_r[144]), .q(net_w[8]));
LSmitll_DFFT_v2p1_optimized DFF_53 (.a(net_r[49]), .clk(net_r[145]), .q(net_w[48]));
LSmitll_DFFT_v2p1_optimized DFF_54 (.a(net_r[50]), .clk(net_r[135]), .q(net_w[49]));
LSmitll_DFFT_v2p1_optimized DFF_55 (.a(net_r[51]), .clk(net_r[134]), .q(net_w[50]));
LSmitll_DFFT_v2p1_optimized DFF_56 (.a(net_r[52]), .clk(net_r[121]), .q(net_w[51]));
LSmitll_DFFT_v2p1_optimized DFF_57 (.a(net_r[53]), .clk(net_r[120]), .q(net_w[52]));
LSmitll_DFFT_v2p1_optimized DFF_58 (.a(net_r[54]), .clk(net_r[122]), .q(net_w[9]));
LSmitll_DFFT_v2p1_optimized DFF_59 (.a(net_r[55]), .clk(net_r[124]), .q(net_w[11]));
LSmitll_DFFT_v2p1_optimized DFF_60 (.a(net_r[56]), .clk(net_r[140]), .q(net_w[15]));
LSmitll_DFFT_v2p1_optimized DFF_61 (.a(net_r[57]), .clk(net_r[153]), .q(net_w[19]));
LSmitll_DFFT_v2p1_optimized DFF_62 (.a(net_r[58]), .clk(net_r[161]), .q(net_w[23]));
LSmitll_DFFT_v2p1_optimized DFF_63 (.a(net_r[59]), .clk(net_r[162]), .q(net_w[25]));
LSmitll_DFFT_v2p1_optimized DFF_64 (.a(net_r[60]), .clk(net_r[156]), .q(net_w[59]));
LSmitll_DFFT_v2p1_optimized DFF_65 (.a(net_r[61]), .clk(net_r[155]), .q(net_w[60]));
LSmitll_DFFT_v2p1_optimized DFF_66 (.a(net_r[62]), .clk(net_r[147]), .q(net_w[61]));
LSmitll_DFFT_v2p1_optimized DFF_67 (.a(net_r[63]), .clk(net_r[146]), .q(net_w[62]));
LSmitll_DFFT_v2p1_optimized DFF_68 (.a(net_r[64]), .clk(net_r[137]), .q(net_w[63]));
LSmitll_DFFT_v2p1_optimized DFF_69 (.a(net_r[65]), .clk(net_r[136]), .q(net_w[64]));
LSmitll_DFFT_v2p1_optimized DFF_70 (.a(net_r[66]), .clk(net_r[163]), .q(net_w[26]));
LSmitll_DFFT_v2p1_optimized DFF_71 (.a(net_r[67]), .clk(net_r[164]), .q(net_w[66]));
LSmitll_DFFT_v2p1_optimized DFF_72 (.a(net_r[68]), .clk(net_r[158]), .q(net_w[67]));
LSmitll_DFFT_v2p1_optimized DFF_73 (.a(net_r[69]), .clk(net_r[157]), .q(net_w[68]));
LSmitll_DFFT_v2p1_optimized DFF_74 (.a(net_r[70]), .clk(net_r[149]), .q(net_w[69]));
LSmitll_DFFT_v2p1_optimized DFF_75 (.a(net_r[71]), .clk(net_r[168]), .q(net_w[27]));
LSmitll_DFFT_v2p1_optimized DFF_76 (.a(net_r[72]), .clk(net_r[165]), .q(net_w[71]));
LSmitll_DFFT_v2p1_optimized DFF_77 (.a(net_r[73]), .clk(net_r[166]), .q(net_w[72]));
LSmitll_DFFT_v2p1_optimized DFF_78 (.a(net_r[74]), .clk(net_r[169]), .q(net_w[28]));
LSmitll_SPLITT_v2p1_optimized SPLIT_79 (.a(net_r[1]), .q(net_w[75]), .m(net_w[76]));
LSmitll_SPLITT_v2p1_optimized SPLIT_80 (.a(net_r[2]), .q(net_w[77]), .m(net_w[78]));
LSmitll_SPLITT_v2p1_optimized SPLIT_81 (.a(net_r[3]), .q(net_w[79]), .m(net_w[80]));
LSmitll_SPLITT_v2p1_optimized SPLIT_82 (.a(net_r[4]), .q(net_w[81]), .m(net_w[82]));
LSmitll_SPLITT_v2p1_optimized SPLIT_83 (.a(net_r[5]), .q(net_w[83]), .m(net_w[84]));
LSmitll_SPLITT_v2p1_optimized SPLIT_84 (.a(net_r[6]), .q(net_w[85]), .m(net_w[86]));
LSmitll_SPLITT_v2p1_optimized SPLIT_85 (.a(net_r[7]), .q(net_w[87]), .m(net_w[88]));
LSmitll_SPLITT_v2p1_optimized SPLIT_86 (.a(net_r[8]), .q(net_w[89]), .m(net_w[90]));
LSmitll_SPLITT_v2p1_optimized SPLIT_87 (.a(net_r[9]), .q(net_w[91]), .m(net_w[92]));
LSmitll_SPLITT_v2p1_optimized SPLIT_88 (.a(net_r[10]), .q(net_w[93]), .m(net_w[94]));
LSmitll_SPLITT_v2p1_optimized SPLIT_89 (.a(net_r[13]), .q(net_w[95]), .m(net_w[96]));
LSmitll_SPLITT_v2p1_optimized SPLIT_90 (.a(net_r[14]), .q(net_w[97]), .m(net_w[98]));
LSmitll_SPLITT_v2p1_optimized SPLIT_91 (.a(net_r[17]), .q(net_w[99]), .m(net_w[100]));
LSmitll_SPLITT_v2p1_optimized SPLIT_92 (.a(net_r[18]), .q(net_w[101]), .m(net_w[102]));
LSmitll_SPLITT_v2p1_optimized SPLIT_93 (.a(net_r[21]), .q(net_w[103]), .m(net_w[104]));
LSmitll_SPLITT_v2p1_optimized SPLIT_94 (.a(net_r[22]), .q(net_w[105]), .m(net_w[106]));
LSmitll_SPLITT_v2p1_optimized SC_96 (.a(net_r[173]), .q(net_w[108]), .m(net_w[109]));
LSmitll_SPLITT_v2p1_optimized SC_97 (.a(net_r[174]), .q(net_w[110]), .m(net_w[111]));
LSmitll_SPLITT_v2p1_optimized SC_98 (.a(net_r[175]), .q(net_w[112]), .m(net_w[113]));
LSmitll_SPLITT_v2p1_optimized SC_99 (.a(net_r[176]), .q(net_w[114]), .m(net_w[115]));
LSmitll_SPLITT_v2p1_optimized SC_100 (.a(net_r[177]), .q(net_w[116]), .m(net_w[117]));
LSmitll_SPLITT_v2p1_optimized SC_101 (.a(net_r[178]), .q(net_w[118]), .m(net_w[119]));
LSmitll_SPLITT_v2p1_optimized SC_102 (.a(net_r[179]), .q(net_w[120]), .m(net_w[121]));
LSmitll_SPLITT_v2p1_optimized SC_103 (.a(net_r[180]), .q(net_w[122]), .m());
LSmitll_SPLITT_v2p1_optimized SC_104 (.a(net_r[187]), .q(net_w[123]), .m(net_w[124]));
LSmitll_SPLITT_v2p1_optimized SC_105 (.a(net_r[188]), .q(net_w[125]), .m(net_w[126]));
LSmitll_SPLITT_v2p1_optimized SC_106 (.a(net_r[189]), .q(net_w[127]), .m(net_w[128]));
LSmitll_SPLITT_v2p1_optimized SC_107 (.a(net_r[190]), .q(net_w[129]), .m(net_w[130]));
LSmitll_SPLITT_v2p1_optimized SC_108 (.a(net_r[191]), .q(net_w[131]), .m(net_w[132]));
LSmitll_SPLITT_v2p1_optimized SC_109 (.a(net_r[192]), .q(net_w[133]), .m(net_w[134]));
LSmitll_SPLITT_v2p1_optimized SC_110 (.a(net_r[193]), .q(net_w[135]), .m());
LSmitll_SPLITT_v2p1_optimized SC_111 (.a(net_r[200]), .q(net_w[136]), .m(net_w[137]));
LSmitll_SPLITT_v2p1_optimized SC_112 (.a(net_r[201]), .q(net_w[138]), .m(net_w[139]));
LSmitll_SPLITT_v2p1_optimized SC_113 (.a(net_r[202]), .q(net_w[140]), .m(net_w[141]));
LSmitll_SPLITT_v2p1_optimized SC_114 (.a(net_r[203]), .q(net_w[142]), .m(net_w[143]));
LSmitll_SPLITT_v2p1_optimized SC_115 (.a(net_r[204]), .q(net_w[144]), .m(net_w[145]));
LSmitll_SPLITT_v2p1_optimized SC_116 (.a(net_r[210]), .q(net_w[146]), .m(net_w[147]));
LSmitll_SPLITT_v2p1_optimized SC_117 (.a(net_r[211]), .q(net_w[148]), .m(net_w[149]));
LSmitll_SPLITT_v2p1_optimized SC_118 (.a(net_r[212]), .q(net_w[150]), .m(net_w[151]));
LSmitll_SPLITT_v2p1_optimized SC_119 (.a(net_r[213]), .q(net_w[152]), .m(net_w[153]));
LSmitll_SPLITT_v2p1_optimized SC_120 (.a(net_r[214]), .q(net_w[154]), .m());
LSmitll_SPLITT_v2p1_optimized SC_121 (.a(net_r[220]), .q(net_w[155]), .m(net_w[156]));
LSmitll_SPLITT_v2p1_optimized SC_122 (.a(net_r[221]), .q(net_w[157]), .m(net_w[158]));
LSmitll_SPLITT_v2p1_optimized SC_123 (.a(net_r[222]), .q(net_w[159]), .m(net_w[160]));
LSmitll_SPLITT_v2p1_optimized SC_124 (.a(net_r[223]), .q(net_w[161]), .m());
LSmitll_SPLITT_v2p1_optimized SC_125 (.a(net_r[227]), .q(net_w[162]), .m(net_w[163]));
LSmitll_SPLITT_v2p1_optimized SC_126 (.a(net_r[228]), .q(net_w[164]), .m(net_w[165]));
LSmitll_SPLITT_v2p1_optimized SC_127 (.a(net_r[229]), .q(net_w[166]), .m(net_w[167]));
LSmitll_SPLITT_v2p1_optimized SC_128 (.a(net_r[233]), .q(net_w[168]), .m(net_w[169]));
LSmitll_SPLITT_v2p1_optimized SC_129 (.a(net_r[234]), .q(net_w[170]), .m(net_w[171]));
LSmitll_SPLITT_v2p1_optimized SC_130 (.a(net_r[235]), .q(net_w[172]), .m());
LSmitll_SPLITT_v2p1_optimized SC_131 (.a(net_r[181]), .q(net_w[173]), .m(net_w[174]));
LSmitll_SPLITT_v2p1_optimized SC_132 (.a(net_r[182]), .q(net_w[175]), .m(net_w[176]));
LSmitll_SPLITT_v2p1_optimized SC_133 (.a(net_r[183]), .q(net_w[177]), .m(net_w[178]));
LSmitll_SPLITT_v2p1_optimized SC_134 (.a(net_r[184]), .q(net_w[179]), .m(net_w[180]));
LSmitll_SPLITT_v2p1_optimized SC_135 (.a(net_r[185]), .q(net_w[181]), .m(net_w[182]));
LSmitll_SPLITT_v2p1_optimized SC_136 (.a(net_r[186]), .q(net_w[183]), .m(net_w[184]));
LSmitll_SPLITT_v2p1_optimized SC_137 (.a(net_r[245]), .q(net_w[185]), .m(net_w[186]));
LSmitll_SPLITT_v2p1_optimized SC_138 (.a(net_r[194]), .q(net_w[187]), .m(net_w[188]));
LSmitll_SPLITT_v2p1_optimized SC_139 (.a(net_r[195]), .q(net_w[189]), .m(net_w[190]));
LSmitll_SPLITT_v2p1_optimized SC_140 (.a(net_r[197]), .q(net_w[191]), .m(net_w[192]));
LSmitll_SPLITT_v2p1_optimized SC_141 (.a(net_r[196]), .q(net_w[193]), .m());
LSmitll_SPLITT_v2p1_optimized SC_142 (.a(net_r[198]), .q(net_w[194]), .m(net_w[195]));
LSmitll_SPLITT_v2p1_optimized SC_143 (.a(net_r[199]), .q(net_w[196]), .m(net_w[197]));
LSmitll_SPLITT_v2p1_optimized SC_144 (.a(net_r[246]), .q(net_w[198]), .m(net_w[199]));
LSmitll_SPLITT_v2p1_optimized SC_145 (.a(net_r[205]), .q(net_w[200]), .m(net_w[201]));
LSmitll_SPLITT_v2p1_optimized SC_146 (.a(net_r[206]), .q(net_w[202]), .m(net_w[203]));
LSmitll_SPLITT_v2p1_optimized SC_147 (.a(net_r[207]), .q(net_w[204]), .m());
LSmitll_SPLITT_v2p1_optimized SC_148 (.a(net_r[208]), .q(net_w[205]), .m(net_w[206]));
LSmitll_SPLITT_v2p1_optimized SC_149 (.a(net_r[209]), .q(net_w[207]), .m());
LSmitll_SPLITT_v2p1_optimized SC_150 (.a(net_r[247]), .q(net_w[208]), .m(net_w[209]));
LSmitll_SPLITT_v2p1_optimized SC_151 (.a(net_r[215]), .q(net_w[210]), .m(net_w[211]));
LSmitll_SPLITT_v2p1_optimized SC_152 (.a(net_r[216]), .q(net_w[212]), .m(net_w[213]));
LSmitll_SPLITT_v2p1_optimized SC_153 (.a(net_r[217]), .q(net_w[214]), .m());
LSmitll_SPLITT_v2p1_optimized SC_154 (.a(net_r[218]), .q(net_w[215]), .m(net_w[216]));
LSmitll_SPLITT_v2p1_optimized SC_155 (.a(net_r[219]), .q(net_w[217]), .m());
LSmitll_SPLITT_v2p1_optimized SC_156 (.a(net_r[248]), .q(net_w[218]), .m(net_w[219]));
LSmitll_SPLITT_v2p1_optimized SC_157 (.a(net_r[224]), .q(net_w[220]), .m(net_w[221]));
LSmitll_SPLITT_v2p1_optimized SC_158 (.a(net_r[225]), .q(net_w[222]), .m(net_w[223]));
LSmitll_SPLITT_v2p1_optimized SC_159 (.a(net_r[226]), .q(net_w[224]), .m(net_w[225]));
LSmitll_SPLITT_v2p1_optimized SC_160 (.a(net_r[249]), .q(net_w[226]), .m());
LSmitll_SPLITT_v2p1_optimized SC_161 (.a(net_r[230]), .q(net_w[227]), .m(net_w[228]));
LSmitll_SPLITT_v2p1_optimized SC_162 (.a(net_r[231]), .q(net_w[229]), .m());
LSmitll_SPLITT_v2p1_optimized SC_163 (.a(net_r[232]), .q(net_w[230]), .m(net_w[231]));
LSmitll_SPLITT_v2p1_optimized SC_164 (.a(net_r[250]), .q(net_w[232]), .m());
LSmitll_SPLITT_v2p1_optimized SC_165 (.a(net_r[236]), .q(net_w[233]), .m(net_w[234]));
LSmitll_SPLITT_v2p1_optimized SC_166 (.a(net_r[237]), .q(net_w[235]), .m());
LSmitll_SPLITT_v2p1_optimized SC_167 (.a(net_r[238]), .q(net_w[236]), .m(net_w[237]));
LSmitll_SPLITT_v2p1_optimized SC_168 (.a(net_r[251]), .q(net_w[238]), .m());
LSmitll_SPLITT_v2p1_optimized SC_169 (.a(net_r[107]), .q(net_w[239]), .m(net_w[240]));
LSmitll_SPLITT_v2p1_optimized SC_170 (.a(net_r[239]), .q(net_w[241]), .m(net_w[242]));
LSmitll_SPLITT_v2p1_optimized SC_171 (.a(net_r[240]), .q(net_w[243]), .m(net_w[244]));
LSmitll_SPLITT_v2p1_optimized SC_172 (.a(net_r[241]), .q(net_w[245]), .m(net_w[246]));
LSmitll_SPLITT_v2p1_optimized SC_173 (.a(net_r[242]), .q(net_w[247]), .m(net_w[248]));
LSmitll_SPLITT_v2p1_optimized SC_174 (.a(net_r[243]), .q(net_w[249]), .m(net_w[250]));
LSmitll_SPLITT_v2p1_optimized SC_175 (.a(net_r[244]), .q(net_w[251]), .m());
endmodule